module axi_clock_converter (
    input wire BUS_CLK ,
    input wire BUS_RSTN,

    //MASTER 0 以太网主机                       MASTER 1 主机                               MASTER 2 主机                               MASTER 3 主机
    output wire [ 1:0] M0_BUS_WR_ADDR_ID   ,    output wire [ 1:0] M1_BUS_WR_ADDR_ID   ,    output wire [ 1:0] M2_BUS_WR_ADDR_ID   ,    output wire [ 1:0] M3_BUS_WR_ADDR_ID   ,
    output wire [31:0] M0_BUS_WR_ADDR      ,    output wire [31:0] M1_BUS_WR_ADDR      ,    output wire [31:0] M2_BUS_WR_ADDR      ,    output wire [31:0] M3_BUS_WR_ADDR      ,
    output wire [ 7:0] M0_BUS_WR_ADDR_LEN  ,    output wire [ 7:0] M1_BUS_WR_ADDR_LEN  ,    output wire [ 7:0] M2_BUS_WR_ADDR_LEN  ,    output wire [ 7:0] M3_BUS_WR_ADDR_LEN  ,
    output wire [ 1:0] M0_BUS_WR_ADDR_BURST,    output wire [ 1:0] M1_BUS_WR_ADDR_BURST,    output wire [ 1:0] M2_BUS_WR_ADDR_BURST,    output wire [ 1:0] M3_BUS_WR_ADDR_BURST,
    output wire        M0_BUS_WR_ADDR_VALID,    output wire        M1_BUS_WR_ADDR_VALID,    output wire        M2_BUS_WR_ADDR_VALID,    output wire        M3_BUS_WR_ADDR_VALID,
    input  wire        M0_BUS_WR_ADDR_READY,    input  wire        M1_BUS_WR_ADDR_READY,    input  wire        M2_BUS_WR_ADDR_READY,    input  wire        M3_BUS_WR_ADDR_READY,

    output wire [31:0] M0_BUS_WR_DATA      ,    output wire [31:0] M1_BUS_WR_DATA      ,    output wire [31:0] M2_BUS_WR_DATA      ,    output wire [31:0] M3_BUS_WR_DATA      ,
    output wire [ 3:0] M0_BUS_WR_STRB      ,    output wire [ 3:0] M1_BUS_WR_STRB      ,    output wire [ 3:0] M2_BUS_WR_STRB      ,    output wire [ 3:0] M3_BUS_WR_STRB      ,
    output wire        M0_BUS_WR_DATA_LAST ,    output wire        M1_BUS_WR_DATA_LAST ,    output wire        M2_BUS_WR_DATA_LAST ,    output wire        M3_BUS_WR_DATA_LAST ,
    output wire        M0_BUS_WR_DATA_VALID,    output wire        M1_BUS_WR_DATA_VALID,    output wire        M2_BUS_WR_DATA_VALID,    output wire        M3_BUS_WR_DATA_VALID,
    input  wire        M0_BUS_WR_DATA_READY,    input  wire        M1_BUS_WR_DATA_READY,    input  wire        M2_BUS_WR_DATA_READY,    input  wire        M3_BUS_WR_DATA_READY,

    input  wire [ 1:0] M0_BUS_WR_BACK_ID   ,    input  wire [ 1:0] M1_BUS_WR_BACK_ID   ,    input  wire [ 1:0] M2_BUS_WR_BACK_ID   ,    input  wire [ 1:0] M3_BUS_WR_BACK_ID   ,
    input  wire [ 1:0] M0_BUS_WR_BACK_RESP ,    input  wire [ 1:0] M1_BUS_WR_BACK_RESP ,    input  wire [ 1:0] M2_BUS_WR_BACK_RESP ,    input  wire [ 1:0] M3_BUS_WR_BACK_RESP ,
    input  wire        M0_BUS_WR_BACK_VALID,    input  wire        M1_BUS_WR_BACK_VALID,    input  wire        M2_BUS_WR_BACK_VALID,    input  wire        M3_BUS_WR_BACK_VALID,
    output wire        M0_BUS_WR_BACK_READY,    output wire        M1_BUS_WR_BACK_READY,    output wire        M2_BUS_WR_BACK_READY,    output wire        M3_BUS_WR_BACK_READY,

    output wire [ 1:0] M0_BUS_RD_ADDR_ID   ,    output wire [ 1:0] M1_BUS_RD_ADDR_ID   ,    output wire [ 1:0] M2_BUS_RD_ADDR_ID   ,    output wire [ 1:0] M3_BUS_RD_ADDR_ID   ,
    output wire [31:0] M0_BUS_RD_ADDR      ,    output wire [31:0] M1_BUS_RD_ADDR      ,    output wire [31:0] M2_BUS_RD_ADDR      ,    output wire [31:0] M3_BUS_RD_ADDR      ,
    output wire [ 7:0] M0_BUS_RD_ADDR_LEN  ,    output wire [ 7:0] M1_BUS_RD_ADDR_LEN  ,    output wire [ 7:0] M2_BUS_RD_ADDR_LEN  ,    output wire [ 7:0] M3_BUS_RD_ADDR_LEN  ,
    output wire [ 1:0] M0_BUS_RD_ADDR_BURST,    output wire [ 1:0] M1_BUS_RD_ADDR_BURST,    output wire [ 1:0] M2_BUS_RD_ADDR_BURST,    output wire [ 1:0] M3_BUS_RD_ADDR_BURST,
    output wire        M0_BUS_RD_ADDR_VALID,    output wire        M1_BUS_RD_ADDR_VALID,    output wire        M2_BUS_RD_ADDR_VALID,    output wire        M3_BUS_RD_ADDR_VALID,
    input  wire        M0_BUS_RD_ADDR_READY,    input  wire        M1_BUS_RD_ADDR_READY,    input  wire        M2_BUS_RD_ADDR_READY,    input  wire        M3_BUS_RD_ADDR_READY,

    input  wire [ 1:0] M0_BUS_RD_BACK_ID   ,    input  wire [ 1:0] M1_BUS_RD_BACK_ID   ,    input  wire [ 1:0] M2_BUS_RD_BACK_ID   ,    input  wire [ 1:0] M3_BUS_RD_BACK_ID   ,
    input  wire [31:0] M0_BUS_RD_DATA      ,    input  wire [31:0] M1_BUS_RD_DATA      ,    input  wire [31:0] M2_BUS_RD_DATA      ,    input  wire [31:0] M3_BUS_RD_DATA      ,
    input  wire [ 1:0] M0_BUS_RD_DATA_RESP ,    input  wire [ 1:0] M1_BUS_RD_DATA_RESP ,    input  wire [ 1:0] M2_BUS_RD_DATA_RESP ,    input  wire [ 1:0] M3_BUS_RD_DATA_RESP ,
    input  wire        M0_BUS_RD_DATA_LAST ,    input  wire        M1_BUS_RD_DATA_LAST ,    input  wire        M2_BUS_RD_DATA_LAST ,    input  wire        M3_BUS_RD_DATA_LAST ,
    input  wire        M0_BUS_RD_DATA_VALID,    input  wire        M1_BUS_RD_DATA_VALID,    input  wire        M2_BUS_RD_DATA_VALID,    input  wire        M3_BUS_RD_DATA_VALID,
    output wire        M0_BUS_RD_DATA_READY,    output wire        M1_BUS_RD_DATA_READY,    output wire        M2_BUS_RD_DATA_READY,    output wire        M3_BUS_RD_DATA_READY,

    //SLAVE 0 DDR从机                           //SLAVE 1 JTAG从机                          //SLAVE 2 从机                              //SLAVE 3 从机
    input  wire [ 3:0] S0_BUS_WR_ADDR_ID   ,    input  wire [ 3:0] S1_BUS_WR_ADDR_ID   ,    input  wire [ 3:0] S2_BUS_WR_ADDR_ID   ,    input  wire [ 3:0] S3_BUS_WR_ADDR_ID   ,
    input  wire [31:0] S0_BUS_WR_ADDR      ,    input  wire [31:0] S1_BUS_WR_ADDR      ,    input  wire [31:0] S2_BUS_WR_ADDR      ,    input  wire [31:0] S3_BUS_WR_ADDR      ,
    input  wire [ 7:0] S0_BUS_WR_ADDR_LEN  ,    input  wire [ 7:0] S1_BUS_WR_ADDR_LEN  ,    input  wire [ 7:0] S2_BUS_WR_ADDR_LEN  ,    input  wire [ 7:0] S3_BUS_WR_ADDR_LEN  ,
    input  wire [ 1:0] S0_BUS_WR_ADDR_BURST,    input  wire [ 1:0] S1_BUS_WR_ADDR_BURST,    input  wire [ 1:0] S2_BUS_WR_ADDR_BURST,    input  wire [ 1:0] S3_BUS_WR_ADDR_BURST,
    input  wire        S0_BUS_WR_ADDR_VALID,    input  wire        S1_BUS_WR_ADDR_VALID,    input  wire        S2_BUS_WR_ADDR_VALID,    input  wire        S3_BUS_WR_ADDR_VALID,
    output wire        S0_BUS_WR_ADDR_READY,    output wire        S1_BUS_WR_ADDR_READY,    output wire        S2_BUS_WR_ADDR_READY,    output wire        S3_BUS_WR_ADDR_READY,

    input  wire [31:0] S0_BUS_WR_DATA      ,    input  wire [31:0] S1_BUS_WR_DATA      ,    input  wire [31:0] S2_BUS_WR_DATA      ,    input  wire [31:0] S3_BUS_WR_DATA      ,
    input  wire [ 3:0] S0_BUS_WR_STRB      ,    input  wire [ 3:0] S1_BUS_WR_STRB      ,    input  wire [ 3:0] S2_BUS_WR_STRB      ,    input  wire [ 3:0] S3_BUS_WR_STRB      ,
    input  wire        S0_BUS_WR_DATA_LAST ,    input  wire        S1_BUS_WR_DATA_LAST ,    input  wire        S2_BUS_WR_DATA_LAST ,    input  wire        S3_BUS_WR_DATA_LAST ,
    input  wire        S0_BUS_WR_DATA_VALID,    input  wire        S1_BUS_WR_DATA_VALID,    input  wire        S2_BUS_WR_DATA_VALID,    input  wire        S3_BUS_WR_DATA_VALID,
    output wire        S0_BUS_WR_DATA_READY,    output wire        S1_BUS_WR_DATA_READY,    output wire        S2_BUS_WR_DATA_READY,    output wire        S3_BUS_WR_DATA_READY,

    output wire [ 3:0] S0_BUS_WR_BACK_ID   ,    output wire [ 3:0] S1_BUS_WR_BACK_ID   ,    output wire [ 3:0] S2_BUS_WR_BACK_ID   ,    output wire [ 3:0] S3_BUS_WR_BACK_ID   ,
    output wire [ 1:0] S0_BUS_WR_BACK_RESP ,    output wire [ 1:0] S1_BUS_WR_BACK_RESP ,    output wire [ 1:0] S2_BUS_WR_BACK_RESP ,    output wire [ 1:0] S3_BUS_WR_BACK_RESP ,
    output wire        S0_BUS_WR_BACK_VALID,    output wire        S1_BUS_WR_BACK_VALID,    output wire        S2_BUS_WR_BACK_VALID,    output wire        S3_BUS_WR_BACK_VALID,
    input  wire        S0_BUS_WR_BACK_READY,    input  wire        S1_BUS_WR_BACK_READY,    input  wire        S2_BUS_WR_BACK_READY,    input  wire        S3_BUS_WR_BACK_READY,

    input  wire [ 3:0] S0_BUS_RD_ADDR_ID   ,    input  wire [ 3:0] S1_BUS_RD_ADDR_ID   ,    input  wire [ 3:0] S2_BUS_RD_ADDR_ID   ,    input  wire [ 3:0] S3_BUS_RD_ADDR_ID   ,
    input  wire [31:0] S0_BUS_RD_ADDR      ,    input  wire [31:0] S1_BUS_RD_ADDR      ,    input  wire [31:0] S2_BUS_RD_ADDR      ,    input  wire [31:0] S3_BUS_RD_ADDR      ,
    input  wire [ 7:0] S0_BUS_RD_ADDR_LEN  ,    input  wire [ 7:0] S1_BUS_RD_ADDR_LEN  ,    input  wire [ 7:0] S2_BUS_RD_ADDR_LEN  ,    input  wire [ 7:0] S3_BUS_RD_ADDR_LEN  ,
    input  wire [ 1:0] S0_BUS_RD_ADDR_BURST,    input  wire [ 1:0] S1_BUS_RD_ADDR_BURST,    input  wire [ 1:0] S2_BUS_RD_ADDR_BURST,    input  wire [ 1:0] S3_BUS_RD_ADDR_BURST,
    input  wire        S0_BUS_RD_ADDR_VALID,    input  wire        S1_BUS_RD_ADDR_VALID,    input  wire        S2_BUS_RD_ADDR_VALID,    input  wire        S3_BUS_RD_ADDR_VALID,
    output wire        S0_BUS_RD_ADDR_READY,    output wire        S1_BUS_RD_ADDR_READY,    output wire        S2_BUS_RD_ADDR_READY,    output wire        S3_BUS_RD_ADDR_READY,

    output wire [ 3:0] S0_BUS_RD_BACK_ID   ,    output wire [ 3:0] S1_BUS_RD_BACK_ID   ,    output wire [ 3:0] S2_BUS_RD_BACK_ID   ,    output wire [ 3:0] S3_BUS_RD_BACK_ID   ,
    output wire [31:0] S0_BUS_RD_DATA      ,    output wire [31:0] S1_BUS_RD_DATA      ,    output wire [31:0] S2_BUS_RD_DATA      ,    output wire [31:0] S3_BUS_RD_DATA      ,
    output wire [ 1:0] S0_BUS_RD_DATA_RESP ,    output wire [ 1:0] S1_BUS_RD_DATA_RESP ,    output wire [ 1:0] S2_BUS_RD_DATA_RESP ,    output wire [ 1:0] S3_BUS_RD_DATA_RESP ,
    output wire        S0_BUS_RD_DATA_LAST ,    output wire        S1_BUS_RD_DATA_LAST ,    output wire        S2_BUS_RD_DATA_LAST ,    output wire        S3_BUS_RD_DATA_LAST ,
    output wire        S0_BUS_RD_DATA_VALID,    output wire        S1_BUS_RD_DATA_VALID,    output wire        S2_BUS_RD_DATA_VALID,    output wire        S3_BUS_RD_DATA_VALID,
    input  wire        S0_BUS_RD_DATA_READY,    input  wire        S1_BUS_RD_DATA_READY,    input  wire        S2_BUS_RD_DATA_READY,    input  wire        S3_BUS_RD_DATA_READY,

    //_______________________________________________________________________________________________________________________________________________________//

    //MASTER 0 以太网主机                   MASTER 1 主机                           MASTER 2 主机                           MASTER 3 主机
    input  wire        M0_CLK          ,    input  wire        M1_CLK          ,    input  wire        M2_CLK          ,    input  wire        M3_CLK          ,
    input  wire        M0_RSTN         ,    input  wire        M1_RSTN         ,    input  wire        M2_RSTN         ,    input  wire        M3_RSTN         ,
    input  wire [ 1:0] M0_WR_ADDR_ID   ,    input  wire [ 1:0] M1_WR_ADDR_ID   ,    input  wire [ 1:0] M2_WR_ADDR_ID   ,    input  wire [ 1:0] M3_WR_ADDR_ID   ,
    input  wire [31:0] M0_WR_ADDR      ,    input  wire [31:0] M1_WR_ADDR      ,    input  wire [31:0] M2_WR_ADDR      ,    input  wire [31:0] M3_WR_ADDR      ,
    input  wire [ 7:0] M0_WR_ADDR_LEN  ,    input  wire [ 7:0] M1_WR_ADDR_LEN  ,    input  wire [ 7:0] M2_WR_ADDR_LEN  ,    input  wire [ 7:0] M3_WR_ADDR_LEN  ,
    input  wire [ 1:0] M0_WR_ADDR_BURST,    input  wire [ 1:0] M1_WR_ADDR_BURST,    input  wire [ 1:0] M2_WR_ADDR_BURST,    input  wire [ 1:0] M3_WR_ADDR_BURST,
    input  wire        M0_WR_ADDR_VALID,    input  wire        M1_WR_ADDR_VALID,    input  wire        M2_WR_ADDR_VALID,    input  wire        M3_WR_ADDR_VALID,
    output wire        M0_WR_ADDR_READY,    output wire        M1_WR_ADDR_READY,    output wire        M2_WR_ADDR_READY,    output wire        M3_WR_ADDR_READY,

    input  wire [31:0] M0_WR_DATA      ,    input  wire [31:0] M1_WR_DATA      ,    input  wire [31:0] M2_WR_DATA      ,    input  wire [31:0] M3_WR_DATA      ,
    input  wire [ 3:0] M0_WR_STRB      ,    input  wire [ 3:0] M1_WR_STRB      ,    input  wire [ 3:0] M2_WR_STRB      ,    input  wire [ 3:0] M3_WR_STRB      ,
    input  wire        M0_WR_DATA_LAST ,    input  wire        M1_WR_DATA_LAST ,    input  wire        M2_WR_DATA_LAST ,    input  wire        M3_WR_DATA_LAST ,
    input  wire        M0_WR_DATA_VALID,    input  wire        M1_WR_DATA_VALID,    input  wire        M2_WR_DATA_VALID,    input  wire        M3_WR_DATA_VALID,
    output wire        M0_WR_DATA_READY,    output wire        M1_WR_DATA_READY,    output wire        M2_WR_DATA_READY,    output wire        M3_WR_DATA_READY,

    output wire [ 1:0] M0_WR_BACK_ID   ,    output wire [ 1:0] M1_WR_BACK_ID   ,    output wire [ 1:0] M2_WR_BACK_ID   ,    output wire [ 1:0] M3_WR_BACK_ID   ,
    output wire [ 1:0] M0_WR_BACK_RESP ,    output wire [ 1:0] M1_WR_BACK_RESP ,    output wire [ 1:0] M2_WR_BACK_RESP ,    output wire [ 1:0] M3_WR_BACK_RESP ,
    output wire        M0_WR_BACK_VALID,    output wire        M1_WR_BACK_VALID,    output wire        M2_WR_BACK_VALID,    output wire        M3_WR_BACK_VALID,
    input  wire        M0_WR_BACK_READY,    input  wire        M1_WR_BACK_READY,    input  wire        M2_WR_BACK_READY,    input  wire        M3_WR_BACK_READY,

    input  wire [ 1:0] M0_RD_ADDR_ID   ,    input  wire [ 1:0] M1_RD_ADDR_ID   ,    input  wire [ 1:0] M2_RD_ADDR_ID   ,    input  wire [ 1:0] M3_RD_ADDR_ID   ,
    input  wire [31:0] M0_RD_ADDR      ,    input  wire [31:0] M1_RD_ADDR      ,    input  wire [31:0] M2_RD_ADDR      ,    input  wire [31:0] M3_RD_ADDR      ,
    input  wire [ 7:0] M0_RD_ADDR_LEN  ,    input  wire [ 7:0] M1_RD_ADDR_LEN  ,    input  wire [ 7:0] M2_RD_ADDR_LEN  ,    input  wire [ 7:0] M3_RD_ADDR_LEN  ,
    input  wire [ 1:0] M0_RD_ADDR_BURST,    input  wire [ 1:0] M1_RD_ADDR_BURST,    input  wire [ 1:0] M2_RD_ADDR_BURST,    input  wire [ 1:0] M3_RD_ADDR_BURST,
    input  wire        M0_RD_ADDR_VALID,    input  wire        M1_RD_ADDR_VALID,    input  wire        M2_RD_ADDR_VALID,    input  wire        M3_RD_ADDR_VALID,
    output wire        M0_RD_ADDR_READY,    output wire        M1_RD_ADDR_READY,    output wire        M2_RD_ADDR_READY,    output wire        M3_RD_ADDR_READY,

    output wire [ 1:0] M0_RD_BACK_ID   ,    output wire [ 1:0] M1_RD_BACK_ID   ,    output wire [ 1:0] M2_RD_BACK_ID   ,    output wire [ 1:0] M3_RD_BACK_ID   ,
    output wire [31:0] M0_RD_DATA      ,    output wire [31:0] M1_RD_DATA      ,    output wire [31:0] M2_RD_DATA      ,    output wire [31:0] M3_RD_DATA      ,
    output wire [ 1:0] M0_RD_DATA_RESP ,    output wire [ 1:0] M1_RD_DATA_RESP ,    output wire [ 1:0] M2_RD_DATA_RESP ,    output wire [ 1:0] M3_RD_DATA_RESP ,
    output wire        M0_RD_DATA_LAST ,    output wire        M1_RD_DATA_LAST ,    output wire        M2_RD_DATA_LAST ,    output wire        M3_RD_DATA_LAST ,
    output wire        M0_RD_DATA_VALID,    output wire        M1_RD_DATA_VALID,    output wire        M2_RD_DATA_VALID,    output wire        M3_RD_DATA_VALID,
    input  wire        M0_RD_DATA_READY,    input  wire        M1_RD_DATA_READY,    input  wire        M2_RD_DATA_READY,    input  wire        M3_RD_DATA_READY,

    //SLAVE 0 DDR从机                       //SLAVE 1 JTAG从机                   //SLAVE 2 从机                  //SLAVE 3 从机
    input  wire        S0_CLK          ,    input  wire        S1_CLK          ,    input  wire        S2_CLK          ,    input  wire        S3_CLK          ,
    input  wire        S0_RSTN         ,    input  wire        S1_RSTN         ,    input  wire        S2_RSTN         ,    input  wire        S3_RSTN         ,
    output wire [ 3:0] S0_WR_ADDR_ID   ,    output wire [ 3:0] S1_WR_ADDR_ID   ,    output wire [ 3:0] S2_WR_ADDR_ID   ,    output wire [ 3:0] S3_WR_ADDR_ID   ,
    output wire [31:0] S0_WR_ADDR      ,    output wire [31:0] S1_WR_ADDR      ,    output wire [31:0] S2_WR_ADDR      ,    output wire [31:0] S3_WR_ADDR      ,
    output wire [ 7:0] S0_WR_ADDR_LEN  ,    output wire [ 7:0] S1_WR_ADDR_LEN  ,    output wire [ 7:0] S2_WR_ADDR_LEN  ,    output wire [ 7:0] S3_WR_ADDR_LEN  ,
    output wire [ 1:0] S0_WR_ADDR_BURST,    output wire [ 1:0] S1_WR_ADDR_BURST,    output wire [ 1:0] S2_WR_ADDR_BURST,    output wire [ 1:0] S3_WR_ADDR_BURST,
    output wire        S0_WR_ADDR_VALID,    output wire        S1_WR_ADDR_VALID,    output wire        S2_WR_ADDR_VALID,    output wire        S3_WR_ADDR_VALID,
    input  wire        S0_WR_ADDR_READY,    input  wire        S1_WR_ADDR_READY,    input  wire        S2_WR_ADDR_READY,    input  wire        S3_WR_ADDR_READY,

    output wire [31:0] S0_WR_DATA      ,    output wire [31:0] S1_WR_DATA      ,    output wire [31:0] S2_WR_DATA      ,    output wire [31:0] S3_WR_DATA      ,
    output wire [ 3:0] S0_WR_STRB      ,    output wire [ 3:0] S1_WR_STRB      ,    output wire [ 3:0] S2_WR_STRB      ,    output wire [ 3:0] S3_WR_STRB      ,
    output wire        S0_WR_DATA_LAST ,    output wire        S1_WR_DATA_LAST ,    output wire        S2_WR_DATA_LAST ,    output wire        S3_WR_DATA_LAST ,
    output wire        S0_WR_DATA_VALID,    output wire        S1_WR_DATA_VALID,    output wire        S2_WR_DATA_VALID,    output wire        S3_WR_DATA_VALID,
    input  wire        S0_WR_DATA_READY,    input  wire        S1_WR_DATA_READY,    input  wire        S2_WR_DATA_READY,    input  wire        S3_WR_DATA_READY,

    input  wire [ 3:0] S0_WR_BACK_ID   ,    input  wire [ 3:0] S1_WR_BACK_ID   ,    input  wire [ 3:0] S2_WR_BACK_ID   ,    input  wire [ 3:0] S3_WR_BACK_ID   ,
    input  wire [ 1:0] S0_WR_BACK_RESP ,    input  wire [ 1:0] S1_WR_BACK_RESP ,    input  wire [ 1:0] S2_WR_BACK_RESP ,    input  wire [ 1:0] S3_WR_BACK_RESP ,
    input  wire        S0_WR_BACK_VALID,    input  wire        S1_WR_BACK_VALID,    input  wire        S2_WR_BACK_VALID,    input  wire        S3_WR_BACK_VALID,
    output wire        S0_WR_BACK_READY,    output wire        S1_WR_BACK_READY,    output wire        S2_WR_BACK_READY,    output wire        S3_WR_BACK_READY,

    output wire [ 3:0] S0_RD_ADDR_ID   ,    output wire [ 3:0] S1_RD_ADDR_ID   ,    output wire [ 3:0] S2_RD_ADDR_ID   ,    output wire [ 3:0] S3_RD_ADDR_ID   ,
    output wire [31:0] S0_RD_ADDR      ,    output wire [31:0] S1_RD_ADDR      ,    output wire [31:0] S2_RD_ADDR      ,    output wire [31:0] S3_RD_ADDR      ,
    output wire [ 7:0] S0_RD_ADDR_LEN  ,    output wire [ 7:0] S1_RD_ADDR_LEN  ,    output wire [ 7:0] S2_RD_ADDR_LEN  ,    output wire [ 7:0] S3_RD_ADDR_LEN  ,
    output wire [ 1:0] S0_RD_ADDR_BURST,    output wire [ 1:0] S1_RD_ADDR_BURST,    output wire [ 1:0] S2_RD_ADDR_BURST,    output wire [ 1:0] S3_RD_ADDR_BURST,
    output wire        S0_RD_ADDR_VALID,    output wire        S1_RD_ADDR_VALID,    output wire        S2_RD_ADDR_VALID,    output wire        S3_RD_ADDR_VALID,
    input  wire        S0_RD_ADDR_READY,    input  wire        S1_RD_ADDR_READY,    input  wire        S2_RD_ADDR_READY,    input  wire        S3_RD_ADDR_READY,

    input  wire [ 3:0] S0_RD_BACK_ID   ,    input  wire [ 3:0] S1_RD_BACK_ID   ,    input  wire [ 3:0] S2_RD_BACK_ID   ,    input  wire [ 3:0] S3_RD_BACK_ID   ,
    input  wire [31:0] S0_RD_DATA      ,    input  wire [31:0] S1_RD_DATA      ,    input  wire [31:0] S2_RD_DATA      ,    input  wire [31:0] S3_RD_DATA      ,
    input  wire [ 1:0] S0_RD_DATA_RESP ,    input  wire [ 1:0] S1_RD_DATA_RESP ,    input  wire [ 1:0] S2_RD_DATA_RESP ,    input  wire [ 1:0] S3_RD_DATA_RESP ,
    input  wire        S0_RD_DATA_LAST ,    input  wire        S1_RD_DATA_LAST ,    input  wire        S2_RD_DATA_LAST ,    input  wire        S3_RD_DATA_LAST ,
    input  wire        S0_RD_DATA_VALID,    input  wire        S1_RD_DATA_VALID,    input  wire        S2_RD_DATA_VALID,    input  wire        S3_RD_DATA_VALID,
    output wire        S0_RD_DATA_READY,    output wire        S1_RD_DATA_READY,    output wire        S2_RD_DATA_READY,    output wire        S3_RD_DATA_READY,
    
    output wire [4:0] M0_fifo_empty_flag, M1_fifo_empty_flag, M2_fifo_empty_flag, M3_fifo_empty_flag,
    output wire [4:0] S0_fifo_empty_flag, S1_fifo_empty_flag, S2_fifo_empty_flag, S3_fifo_empty_flag
);
/*
AXI CLOCK CONVERTER模块，集中处理各个模块的时钟域转换
fifo的引入同时使主从模块支持了outstanding功能
*/

master_axi_async m0_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .MASTER_CLK              (M0_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .MASTER_RSTN             (M0_RSTN         ),
    .BUS_WR_ADDR_ID         (M0_BUS_WR_ADDR_ID   ), /* <===> */ .MASTER_WR_ADDR_ID       (M0_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (M0_BUS_WR_ADDR      ), /* <===> */ .MASTER_WR_ADDR          (M0_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (M0_BUS_WR_ADDR_LEN  ), /* <===> */ .MASTER_WR_ADDR_LEN      (M0_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (M0_BUS_WR_ADDR_BURST), /* <===> */ .MASTER_WR_ADDR_BURST    (M0_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (M0_BUS_WR_ADDR_VALID), /* <===> */ .MASTER_WR_ADDR_VALID    (M0_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (M0_BUS_WR_ADDR_READY), /* <===> */ .MASTER_WR_ADDR_READY    (M0_WR_ADDR_READY),
    .BUS_WR_DATA            (M0_BUS_WR_DATA      ), /* <===> */ .MASTER_WR_DATA          (M0_WR_DATA      ),
    .BUS_WR_STRB            (M0_BUS_WR_STRB      ), /* <===> */ .MASTER_WR_STRB          (M0_WR_STRB      ),
    .BUS_WR_DATA_LAST       (M0_BUS_WR_DATA_LAST ), /* <===> */ .MASTER_WR_DATA_LAST     (M0_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (M0_BUS_WR_DATA_VALID), /* <===> */ .MASTER_WR_DATA_VALID    (M0_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (M0_BUS_WR_DATA_READY), /* <===> */ .MASTER_WR_DATA_READY    (M0_WR_DATA_READY),
    .BUS_WR_BACK_ID         (M0_BUS_WR_BACK_ID   ), /* <===> */ .MASTER_WR_BACK_ID       (M0_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (M0_BUS_WR_BACK_RESP ), /* <===> */ .MASTER_WR_BACK_RESP     (M0_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (M0_BUS_WR_BACK_VALID), /* <===> */ .MASTER_WR_BACK_VALID    (M0_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (M0_BUS_WR_BACK_READY), /* <===> */ .MASTER_WR_BACK_READY    (M0_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (M0_BUS_RD_ADDR_ID   ), /* <===> */ .MASTER_RD_ADDR_ID       (M0_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (M0_BUS_RD_ADDR      ), /* <===> */ .MASTER_RD_ADDR          (M0_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (M0_BUS_RD_ADDR_LEN  ), /* <===> */ .MASTER_RD_ADDR_LEN      (M0_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (M0_BUS_RD_ADDR_BURST), /* <===> */ .MASTER_RD_ADDR_BURST    (M0_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (M0_BUS_RD_ADDR_VALID), /* <===> */ .MASTER_RD_ADDR_VALID    (M0_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (M0_BUS_RD_ADDR_READY), /* <===> */ .MASTER_RD_ADDR_READY    (M0_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (M0_BUS_RD_BACK_ID   ), /* <===> */ .MASTER_RD_BACK_ID       (M0_RD_BACK_ID   ),
    .BUS_RD_DATA            (M0_BUS_RD_DATA      ), /* <===> */ .MASTER_RD_DATA          (M0_RD_DATA      ),
    .BUS_RD_DATA_RESP       (M0_BUS_RD_DATA_RESP ), /* <===> */ .MASTER_RD_DATA_RESP     (M0_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (M0_BUS_RD_DATA_LAST ), /* <===> */ .MASTER_RD_DATA_LAST     (M0_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (M0_BUS_RD_DATA_VALID), /* <===> */ .MASTER_RD_DATA_VALID    (M0_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (M0_BUS_RD_DATA_READY), /* <===> */ .MASTER_RD_DATA_READY    (M0_RD_DATA_READY),
    .fifo_empty_flag        (M0_fifo_empty_flag)
);

master_axi_async m1_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .MASTER_CLK              (M1_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .MASTER_RSTN             (M1_RSTN         ),
    .BUS_WR_ADDR_ID         (M1_BUS_WR_ADDR_ID   ), /* <===> */ .MASTER_WR_ADDR_ID       (M1_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (M1_BUS_WR_ADDR      ), /* <===> */ .MASTER_WR_ADDR          (M1_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (M1_BUS_WR_ADDR_LEN  ), /* <===> */ .MASTER_WR_ADDR_LEN      (M1_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (M1_BUS_WR_ADDR_BURST), /* <===> */ .MASTER_WR_ADDR_BURST    (M1_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (M1_BUS_WR_ADDR_VALID), /* <===> */ .MASTER_WR_ADDR_VALID    (M1_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (M1_BUS_WR_ADDR_READY), /* <===> */ .MASTER_WR_ADDR_READY    (M1_WR_ADDR_READY),
    .BUS_WR_DATA            (M1_BUS_WR_DATA      ), /* <===> */ .MASTER_WR_DATA          (M1_WR_DATA      ),
    .BUS_WR_STRB            (M1_BUS_WR_STRB      ), /* <===> */ .MASTER_WR_STRB          (M1_WR_STRB      ),
    .BUS_WR_DATA_LAST       (M1_BUS_WR_DATA_LAST ), /* <===> */ .MASTER_WR_DATA_LAST     (M1_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (M1_BUS_WR_DATA_VALID), /* <===> */ .MASTER_WR_DATA_VALID    (M1_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (M1_BUS_WR_DATA_READY), /* <===> */ .MASTER_WR_DATA_READY    (M1_WR_DATA_READY),
    .BUS_WR_BACK_ID         (M1_BUS_WR_BACK_ID   ), /* <===> */ .MASTER_WR_BACK_ID       (M1_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (M1_BUS_WR_BACK_RESP ), /* <===> */ .MASTER_WR_BACK_RESP     (M1_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (M1_BUS_WR_BACK_VALID), /* <===> */ .MASTER_WR_BACK_VALID    (M1_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (M1_BUS_WR_BACK_READY), /* <===> */ .MASTER_WR_BACK_READY    (M1_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (M1_BUS_RD_ADDR_ID   ), /* <===> */ .MASTER_RD_ADDR_ID       (M1_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (M1_BUS_RD_ADDR      ), /* <===> */ .MASTER_RD_ADDR          (M1_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (M1_BUS_RD_ADDR_LEN  ), /* <===> */ .MASTER_RD_ADDR_LEN      (M1_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (M1_BUS_RD_ADDR_BURST), /* <===> */ .MASTER_RD_ADDR_BURST    (M1_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (M1_BUS_RD_ADDR_VALID), /* <===> */ .MASTER_RD_ADDR_VALID    (M1_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (M1_BUS_RD_ADDR_READY), /* <===> */ .MASTER_RD_ADDR_READY    (M1_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (M1_BUS_RD_BACK_ID   ), /* <===> */ .MASTER_RD_BACK_ID       (M1_RD_BACK_ID   ),
    .BUS_RD_DATA            (M1_BUS_RD_DATA      ), /* <===> */ .MASTER_RD_DATA          (M1_RD_DATA      ),
    .BUS_RD_DATA_RESP       (M1_BUS_RD_DATA_RESP ), /* <===> */ .MASTER_RD_DATA_RESP     (M1_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (M1_BUS_RD_DATA_LAST ), /* <===> */ .MASTER_RD_DATA_LAST     (M1_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (M1_BUS_RD_DATA_VALID), /* <===> */ .MASTER_RD_DATA_VALID    (M1_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (M1_BUS_RD_DATA_READY), /* <===> */ .MASTER_RD_DATA_READY    (M1_RD_DATA_READY),
    .fifo_empty_flag        (M1_fifo_empty_flag)
);

master_axi_async m2_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .MASTER_CLK              (M2_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .MASTER_RSTN             (M2_RSTN         ),
    .BUS_WR_ADDR_ID         (M2_BUS_WR_ADDR_ID   ), /* <===> */ .MASTER_WR_ADDR_ID       (M2_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (M2_BUS_WR_ADDR      ), /* <===> */ .MASTER_WR_ADDR          (M2_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (M2_BUS_WR_ADDR_LEN  ), /* <===> */ .MASTER_WR_ADDR_LEN      (M2_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (M2_BUS_WR_ADDR_BURST), /* <===> */ .MASTER_WR_ADDR_BURST    (M2_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (M2_BUS_WR_ADDR_VALID), /* <===> */ .MASTER_WR_ADDR_VALID    (M2_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (M2_BUS_WR_ADDR_READY), /* <===> */ .MASTER_WR_ADDR_READY    (M2_WR_ADDR_READY),
    .BUS_WR_DATA            (M2_BUS_WR_DATA      ), /* <===> */ .MASTER_WR_DATA          (M2_WR_DATA      ),
    .BUS_WR_STRB            (M2_BUS_WR_STRB      ), /* <===> */ .MASTER_WR_STRB          (M2_WR_STRB      ),
    .BUS_WR_DATA_LAST       (M2_BUS_WR_DATA_LAST ), /* <===> */ .MASTER_WR_DATA_LAST     (M2_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (M2_BUS_WR_DATA_VALID), /* <===> */ .MASTER_WR_DATA_VALID    (M2_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (M2_BUS_WR_DATA_READY), /* <===> */ .MASTER_WR_DATA_READY    (M2_WR_DATA_READY),
    .BUS_WR_BACK_ID         (M2_BUS_WR_BACK_ID   ), /* <===> */ .MASTER_WR_BACK_ID       (M2_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (M2_BUS_WR_BACK_RESP ), /* <===> */ .MASTER_WR_BACK_RESP     (M2_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (M2_BUS_WR_BACK_VALID), /* <===> */ .MASTER_WR_BACK_VALID    (M2_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (M2_BUS_WR_BACK_READY), /* <===> */ .MASTER_WR_BACK_READY    (M2_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (M2_BUS_RD_ADDR_ID   ), /* <===> */ .MASTER_RD_ADDR_ID       (M2_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (M2_BUS_RD_ADDR      ), /* <===> */ .MASTER_RD_ADDR          (M2_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (M2_BUS_RD_ADDR_LEN  ), /* <===> */ .MASTER_RD_ADDR_LEN      (M2_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (M2_BUS_RD_ADDR_BURST), /* <===> */ .MASTER_RD_ADDR_BURST    (M2_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (M2_BUS_RD_ADDR_VALID), /* <===> */ .MASTER_RD_ADDR_VALID    (M2_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (M2_BUS_RD_ADDR_READY), /* <===> */ .MASTER_RD_ADDR_READY    (M2_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (M2_BUS_RD_BACK_ID   ), /* <===> */ .MASTER_RD_BACK_ID       (M2_RD_BACK_ID   ),
    .BUS_RD_DATA            (M2_BUS_RD_DATA      ), /* <===> */ .MASTER_RD_DATA          (M2_RD_DATA      ),
    .BUS_RD_DATA_RESP       (M2_BUS_RD_DATA_RESP ), /* <===> */ .MASTER_RD_DATA_RESP     (M2_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (M2_BUS_RD_DATA_LAST ), /* <===> */ .MASTER_RD_DATA_LAST     (M2_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (M2_BUS_RD_DATA_VALID), /* <===> */ .MASTER_RD_DATA_VALID    (M2_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (M2_BUS_RD_DATA_READY), /* <===> */ .MASTER_RD_DATA_READY    (M2_RD_DATA_READY),
    .fifo_empty_flag        (M2_fifo_empty_flag)
);

master_axi_async m3_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .MASTER_CLK              (M3_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .MASTER_RSTN             (M3_RSTN         ),
    .BUS_WR_ADDR_ID         (M3_BUS_WR_ADDR_ID   ), /* <===> */ .MASTER_WR_ADDR_ID       (M3_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (M3_BUS_WR_ADDR      ), /* <===> */ .MASTER_WR_ADDR          (M3_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (M3_BUS_WR_ADDR_LEN  ), /* <===> */ .MASTER_WR_ADDR_LEN      (M3_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (M3_BUS_WR_ADDR_BURST), /* <===> */ .MASTER_WR_ADDR_BURST    (M3_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (M3_BUS_WR_ADDR_VALID), /* <===> */ .MASTER_WR_ADDR_VALID    (M3_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (M3_BUS_WR_ADDR_READY), /* <===> */ .MASTER_WR_ADDR_READY    (M3_WR_ADDR_READY),
    .BUS_WR_DATA            (M3_BUS_WR_DATA      ), /* <===> */ .MASTER_WR_DATA          (M3_WR_DATA      ),
    .BUS_WR_STRB            (M3_BUS_WR_STRB      ), /* <===> */ .MASTER_WR_STRB          (M3_WR_STRB      ),
    .BUS_WR_DATA_LAST       (M3_BUS_WR_DATA_LAST ), /* <===> */ .MASTER_WR_DATA_LAST     (M3_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (M3_BUS_WR_DATA_VALID), /* <===> */ .MASTER_WR_DATA_VALID    (M3_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (M3_BUS_WR_DATA_READY), /* <===> */ .MASTER_WR_DATA_READY    (M3_WR_DATA_READY),
    .BUS_WR_BACK_ID         (M3_BUS_WR_BACK_ID   ), /* <===> */ .MASTER_WR_BACK_ID       (M3_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (M3_BUS_WR_BACK_RESP ), /* <===> */ .MASTER_WR_BACK_RESP     (M3_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (M3_BUS_WR_BACK_VALID), /* <===> */ .MASTER_WR_BACK_VALID    (M3_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (M3_BUS_WR_BACK_READY), /* <===> */ .MASTER_WR_BACK_READY    (M3_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (M3_BUS_RD_ADDR_ID   ), /* <===> */ .MASTER_RD_ADDR_ID       (M3_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (M3_BUS_RD_ADDR      ), /* <===> */ .MASTER_RD_ADDR          (M3_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (M3_BUS_RD_ADDR_LEN  ), /* <===> */ .MASTER_RD_ADDR_LEN      (M3_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (M3_BUS_RD_ADDR_BURST), /* <===> */ .MASTER_RD_ADDR_BURST    (M3_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (M3_BUS_RD_ADDR_VALID), /* <===> */ .MASTER_RD_ADDR_VALID    (M3_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (M3_BUS_RD_ADDR_READY), /* <===> */ .MASTER_RD_ADDR_READY    (M3_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (M3_BUS_RD_BACK_ID   ), /* <===> */ .MASTER_RD_BACK_ID       (M3_RD_BACK_ID   ),
    .BUS_RD_DATA            (M3_BUS_RD_DATA      ), /* <===> */ .MASTER_RD_DATA          (M3_RD_DATA      ),
    .BUS_RD_DATA_RESP       (M3_BUS_RD_DATA_RESP ), /* <===> */ .MASTER_RD_DATA_RESP     (M3_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (M3_BUS_RD_DATA_LAST ), /* <===> */ .MASTER_RD_DATA_LAST     (M3_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (M3_BUS_RD_DATA_VALID), /* <===> */ .MASTER_RD_DATA_VALID    (M3_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (M3_BUS_RD_DATA_READY), /* <===> */ .MASTER_RD_DATA_READY    (M3_RD_DATA_READY),
    .fifo_empty_flag        (M3_fifo_empty_flag)
);

slave_axi_async s0_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .SLAVE_CLK              (S0_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .SLAVE_RSTN             (S0_RSTN         ),
    .BUS_WR_ADDR_ID         (S0_BUS_WR_ADDR_ID   ), /* <===> */ .SLAVE_WR_ADDR_ID       (S0_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (S0_BUS_WR_ADDR      ), /* <===> */ .SLAVE_WR_ADDR          (S0_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (S0_BUS_WR_ADDR_LEN  ), /* <===> */ .SLAVE_WR_ADDR_LEN      (S0_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (S0_BUS_WR_ADDR_BURST), /* <===> */ .SLAVE_WR_ADDR_BURST    (S0_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (S0_BUS_WR_ADDR_VALID), /* <===> */ .SLAVE_WR_ADDR_VALID    (S0_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (S0_BUS_WR_ADDR_READY), /* <===> */ .SLAVE_WR_ADDR_READY    (S0_WR_ADDR_READY),
    .BUS_WR_DATA            (S0_BUS_WR_DATA      ), /* <===> */ .SLAVE_WR_DATA          (S0_WR_DATA      ),
    .BUS_WR_STRB            (S0_BUS_WR_STRB      ), /* <===> */ .SLAVE_WR_STRB          (S0_WR_STRB      ),
    .BUS_WR_DATA_LAST       (S0_BUS_WR_DATA_LAST ), /* <===> */ .SLAVE_WR_DATA_LAST     (S0_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (S0_BUS_WR_DATA_VALID), /* <===> */ .SLAVE_WR_DATA_VALID    (S0_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (S0_BUS_WR_DATA_READY), /* <===> */ .SLAVE_WR_DATA_READY    (S0_WR_DATA_READY),
    .BUS_WR_BACK_ID         (S0_BUS_WR_BACK_ID   ), /* <===> */ .SLAVE_WR_BACK_ID       (S0_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (S0_BUS_WR_BACK_RESP ), /* <===> */ .SLAVE_WR_BACK_RESP     (S0_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (S0_BUS_WR_BACK_VALID), /* <===> */ .SLAVE_WR_BACK_VALID    (S0_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (S0_BUS_WR_BACK_READY), /* <===> */ .SLAVE_WR_BACK_READY    (S0_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (S0_BUS_RD_ADDR_ID   ), /* <===> */ .SLAVE_RD_ADDR_ID       (S0_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (S0_BUS_RD_ADDR      ), /* <===> */ .SLAVE_RD_ADDR          (S0_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (S0_BUS_RD_ADDR_LEN  ), /* <===> */ .SLAVE_RD_ADDR_LEN      (S0_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (S0_BUS_RD_ADDR_BURST), /* <===> */ .SLAVE_RD_ADDR_BURST    (S0_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (S0_BUS_RD_ADDR_VALID), /* <===> */ .SLAVE_RD_ADDR_VALID    (S0_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (S0_BUS_RD_ADDR_READY), /* <===> */ .SLAVE_RD_ADDR_READY    (S0_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (S0_BUS_RD_BACK_ID   ), /* <===> */ .SLAVE_RD_BACK_ID       (S0_RD_BACK_ID   ),
    .BUS_RD_DATA            (S0_BUS_RD_DATA      ), /* <===> */ .SLAVE_RD_DATA          (S0_RD_DATA      ),
    .BUS_RD_DATA_RESP       (S0_BUS_RD_DATA_RESP ), /* <===> */ .SLAVE_RD_DATA_RESP     (S0_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (S0_BUS_RD_DATA_LAST ), /* <===> */ .SLAVE_RD_DATA_LAST     (S0_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (S0_BUS_RD_DATA_VALID), /* <===> */ .SLAVE_RD_DATA_VALID    (S0_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (S0_BUS_RD_DATA_READY), /* <===> */ .SLAVE_RD_DATA_READY    (S0_RD_DATA_READY),
    .fifo_empty_flag        (S0_fifo_empty_flag)
);

slave_axi_async s1_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .SLAVE_CLK              (S1_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .SLAVE_RSTN             (S1_RSTN         ),
    .BUS_WR_ADDR_ID         (S1_BUS_WR_ADDR_ID   ), /* <===> */ .SLAVE_WR_ADDR_ID       (S1_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (S1_BUS_WR_ADDR      ), /* <===> */ .SLAVE_WR_ADDR          (S1_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (S1_BUS_WR_ADDR_LEN  ), /* <===> */ .SLAVE_WR_ADDR_LEN      (S1_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (S1_BUS_WR_ADDR_BURST), /* <===> */ .SLAVE_WR_ADDR_BURST    (S1_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (S1_BUS_WR_ADDR_VALID), /* <===> */ .SLAVE_WR_ADDR_VALID    (S1_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (S1_BUS_WR_ADDR_READY), /* <===> */ .SLAVE_WR_ADDR_READY    (S1_WR_ADDR_READY),
    .BUS_WR_DATA            (S1_BUS_WR_DATA      ), /* <===> */ .SLAVE_WR_DATA          (S1_WR_DATA      ),
    .BUS_WR_STRB            (S1_BUS_WR_STRB      ), /* <===> */ .SLAVE_WR_STRB          (S1_WR_STRB      ),
    .BUS_WR_DATA_LAST       (S1_BUS_WR_DATA_LAST ), /* <===> */ .SLAVE_WR_DATA_LAST     (S1_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (S1_BUS_WR_DATA_VALID), /* <===> */ .SLAVE_WR_DATA_VALID    (S1_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (S1_BUS_WR_DATA_READY), /* <===> */ .SLAVE_WR_DATA_READY    (S1_WR_DATA_READY),
    .BUS_WR_BACK_ID         (S1_BUS_WR_BACK_ID   ), /* <===> */ .SLAVE_WR_BACK_ID       (S1_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (S1_BUS_WR_BACK_RESP ), /* <===> */ .SLAVE_WR_BACK_RESP     (S1_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (S1_BUS_WR_BACK_VALID), /* <===> */ .SLAVE_WR_BACK_VALID    (S1_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (S1_BUS_WR_BACK_READY), /* <===> */ .SLAVE_WR_BACK_READY    (S1_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (S1_BUS_RD_ADDR_ID   ), /* <===> */ .SLAVE_RD_ADDR_ID       (S1_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (S1_BUS_RD_ADDR      ), /* <===> */ .SLAVE_RD_ADDR          (S1_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (S1_BUS_RD_ADDR_LEN  ), /* <===> */ .SLAVE_RD_ADDR_LEN      (S1_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (S1_BUS_RD_ADDR_BURST), /* <===> */ .SLAVE_RD_ADDR_BURST    (S1_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (S1_BUS_RD_ADDR_VALID), /* <===> */ .SLAVE_RD_ADDR_VALID    (S1_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (S1_BUS_RD_ADDR_READY), /* <===> */ .SLAVE_RD_ADDR_READY    (S1_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (S1_BUS_RD_BACK_ID   ), /* <===> */ .SLAVE_RD_BACK_ID       (S1_RD_BACK_ID   ),
    .BUS_RD_DATA            (S1_BUS_RD_DATA      ), /* <===> */ .SLAVE_RD_DATA          (S1_RD_DATA      ),
    .BUS_RD_DATA_RESP       (S1_BUS_RD_DATA_RESP ), /* <===> */ .SLAVE_RD_DATA_RESP     (S1_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (S1_BUS_RD_DATA_LAST ), /* <===> */ .SLAVE_RD_DATA_LAST     (S1_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (S1_BUS_RD_DATA_VALID), /* <===> */ .SLAVE_RD_DATA_VALID    (S1_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (S1_BUS_RD_DATA_READY), /* <===> */ .SLAVE_RD_DATA_READY    (S1_RD_DATA_READY),
    .fifo_empty_flag        (S1_fifo_empty_flag)
);

slave_axi_async s2_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .SLAVE_CLK              (S2_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .SLAVE_RSTN             (S2_RSTN         ),
    .BUS_WR_ADDR_ID         (S2_BUS_WR_ADDR_ID   ), /* <===> */ .SLAVE_WR_ADDR_ID       (S2_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (S2_BUS_WR_ADDR      ), /* <===> */ .SLAVE_WR_ADDR          (S2_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (S2_BUS_WR_ADDR_LEN  ), /* <===> */ .SLAVE_WR_ADDR_LEN      (S2_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (S2_BUS_WR_ADDR_BURST), /* <===> */ .SLAVE_WR_ADDR_BURST    (S2_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (S2_BUS_WR_ADDR_VALID), /* <===> */ .SLAVE_WR_ADDR_VALID    (S2_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (S2_BUS_WR_ADDR_READY), /* <===> */ .SLAVE_WR_ADDR_READY    (S2_WR_ADDR_READY),
    .BUS_WR_DATA            (S2_BUS_WR_DATA      ), /* <===> */ .SLAVE_WR_DATA          (S2_WR_DATA      ),
    .BUS_WR_STRB            (S2_BUS_WR_STRB      ), /* <===> */ .SLAVE_WR_STRB          (S2_WR_STRB      ),
    .BUS_WR_DATA_LAST       (S2_BUS_WR_DATA_LAST ), /* <===> */ .SLAVE_WR_DATA_LAST     (S2_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (S2_BUS_WR_DATA_VALID), /* <===> */ .SLAVE_WR_DATA_VALID    (S2_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (S2_BUS_WR_DATA_READY), /* <===> */ .SLAVE_WR_DATA_READY    (S2_WR_DATA_READY),
    .BUS_WR_BACK_ID         (S2_BUS_WR_BACK_ID   ), /* <===> */ .SLAVE_WR_BACK_ID       (S2_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (S2_BUS_WR_BACK_RESP ), /* <===> */ .SLAVE_WR_BACK_RESP     (S2_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (S2_BUS_WR_BACK_VALID), /* <===> */ .SLAVE_WR_BACK_VALID    (S2_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (S2_BUS_WR_BACK_READY), /* <===> */ .SLAVE_WR_BACK_READY    (S2_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (S2_BUS_RD_ADDR_ID   ), /* <===> */ .SLAVE_RD_ADDR_ID       (S2_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (S2_BUS_RD_ADDR      ), /* <===> */ .SLAVE_RD_ADDR          (S2_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (S2_BUS_RD_ADDR_LEN  ), /* <===> */ .SLAVE_RD_ADDR_LEN      (S2_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (S2_BUS_RD_ADDR_BURST), /* <===> */ .SLAVE_RD_ADDR_BURST    (S2_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (S2_BUS_RD_ADDR_VALID), /* <===> */ .SLAVE_RD_ADDR_VALID    (S2_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (S2_BUS_RD_ADDR_READY), /* <===> */ .SLAVE_RD_ADDR_READY    (S2_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (S2_BUS_RD_BACK_ID   ), /* <===> */ .SLAVE_RD_BACK_ID       (S2_RD_BACK_ID   ),
    .BUS_RD_DATA            (S2_BUS_RD_DATA      ), /* <===> */ .SLAVE_RD_DATA          (S2_RD_DATA      ),
    .BUS_RD_DATA_RESP       (S2_BUS_RD_DATA_RESP ), /* <===> */ .SLAVE_RD_DATA_RESP     (S2_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (S2_BUS_RD_DATA_LAST ), /* <===> */ .SLAVE_RD_DATA_LAST     (S2_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (S2_BUS_RD_DATA_VALID), /* <===> */ .SLAVE_RD_DATA_VALID    (S2_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (S2_BUS_RD_DATA_READY), /* <===> */ .SLAVE_RD_DATA_READY    (S2_RD_DATA_READY),
    .fifo_empty_flag        (S2_fifo_empty_flag)
);

slave_axi_async s3_axi_async(
    .BUS_CLK                (   BUS_CLK          ), /* <===> */ .SLAVE_CLK              (S3_CLK          ),
    .BUS_RSTN               (   BUS_RSTN         ), /* <===> */ .SLAVE_RSTN             (S3_RSTN         ),
    .BUS_WR_ADDR_ID         (S3_BUS_WR_ADDR_ID   ), /* <===> */ .SLAVE_WR_ADDR_ID       (S3_WR_ADDR_ID   ),
    .BUS_WR_ADDR            (S3_BUS_WR_ADDR      ), /* <===> */ .SLAVE_WR_ADDR          (S3_WR_ADDR      ),
    .BUS_WR_ADDR_LEN        (S3_BUS_WR_ADDR_LEN  ), /* <===> */ .SLAVE_WR_ADDR_LEN      (S3_WR_ADDR_LEN  ),
    .BUS_WR_ADDR_BURST      (S3_BUS_WR_ADDR_BURST), /* <===> */ .SLAVE_WR_ADDR_BURST    (S3_WR_ADDR_BURST),
    .BUS_WR_ADDR_VALID      (S3_BUS_WR_ADDR_VALID), /* <===> */ .SLAVE_WR_ADDR_VALID    (S3_WR_ADDR_VALID),
    .BUS_WR_ADDR_READY      (S3_BUS_WR_ADDR_READY), /* <===> */ .SLAVE_WR_ADDR_READY    (S3_WR_ADDR_READY),
    .BUS_WR_DATA            (S3_BUS_WR_DATA      ), /* <===> */ .SLAVE_WR_DATA          (S3_WR_DATA      ),
    .BUS_WR_STRB            (S3_BUS_WR_STRB      ), /* <===> */ .SLAVE_WR_STRB          (S3_WR_STRB      ),
    .BUS_WR_DATA_LAST       (S3_BUS_WR_DATA_LAST ), /* <===> */ .SLAVE_WR_DATA_LAST     (S3_WR_DATA_LAST ),
    .BUS_WR_DATA_VALID      (S3_BUS_WR_DATA_VALID), /* <===> */ .SLAVE_WR_DATA_VALID    (S3_WR_DATA_VALID),
    .BUS_WR_DATA_READY      (S3_BUS_WR_DATA_READY), /* <===> */ .SLAVE_WR_DATA_READY    (S3_WR_DATA_READY),
    .BUS_WR_BACK_ID         (S3_BUS_WR_BACK_ID   ), /* <===> */ .SLAVE_WR_BACK_ID       (S3_WR_BACK_ID   ),
    .BUS_WR_BACK_RESP       (S3_BUS_WR_BACK_RESP ), /* <===> */ .SLAVE_WR_BACK_RESP     (S3_WR_BACK_RESP ),
    .BUS_WR_BACK_VALID      (S3_BUS_WR_BACK_VALID), /* <===> */ .SLAVE_WR_BACK_VALID    (S3_WR_BACK_VALID),
    .BUS_WR_BACK_READY      (S3_BUS_WR_BACK_READY), /* <===> */ .SLAVE_WR_BACK_READY    (S3_WR_BACK_READY),
    .BUS_RD_ADDR_ID         (S3_BUS_RD_ADDR_ID   ), /* <===> */ .SLAVE_RD_ADDR_ID       (S3_RD_ADDR_ID   ),
    .BUS_RD_ADDR            (S3_BUS_RD_ADDR      ), /* <===> */ .SLAVE_RD_ADDR          (S3_RD_ADDR      ),
    .BUS_RD_ADDR_LEN        (S3_BUS_RD_ADDR_LEN  ), /* <===> */ .SLAVE_RD_ADDR_LEN      (S3_RD_ADDR_LEN  ),
    .BUS_RD_ADDR_BURST      (S3_BUS_RD_ADDR_BURST), /* <===> */ .SLAVE_RD_ADDR_BURST    (S3_RD_ADDR_BURST),
    .BUS_RD_ADDR_VALID      (S3_BUS_RD_ADDR_VALID), /* <===> */ .SLAVE_RD_ADDR_VALID    (S3_RD_ADDR_VALID),
    .BUS_RD_ADDR_READY      (S3_BUS_RD_ADDR_READY), /* <===> */ .SLAVE_RD_ADDR_READY    (S3_RD_ADDR_READY),
    .BUS_RD_BACK_ID         (S3_BUS_RD_BACK_ID   ), /* <===> */ .SLAVE_RD_BACK_ID       (S3_RD_BACK_ID   ),
    .BUS_RD_DATA            (S3_BUS_RD_DATA      ), /* <===> */ .SLAVE_RD_DATA          (S3_RD_DATA      ),
    .BUS_RD_DATA_RESP       (S3_BUS_RD_DATA_RESP ), /* <===> */ .SLAVE_RD_DATA_RESP     (S3_RD_DATA_RESP ),
    .BUS_RD_DATA_LAST       (S3_BUS_RD_DATA_LAST ), /* <===> */ .SLAVE_RD_DATA_LAST     (S3_RD_DATA_LAST ),
    .BUS_RD_DATA_VALID      (S3_BUS_RD_DATA_VALID), /* <===> */ .SLAVE_RD_DATA_VALID    (S3_RD_DATA_VALID),
    .BUS_RD_DATA_READY      (S3_BUS_RD_DATA_READY), /* <===> */ .SLAVE_RD_DATA_READY    (S3_RD_DATA_READY),
    .fifo_empty_flag        (S3_fifo_empty_flag)
);

endmodule