`timescale 1ns/1ps
module remote_update_test ();

reg BUS_CLK;
reg BUS_RSTN;

localparam M_WIDTH  = 2;
localparam S_WIDTH  = 2;
localparam M_ID     = 2;
localparam [0:(2**S_WIDTH-1)][31:0] START_ADDR = {32'h00000000, 32'h10000000, 32'h20000000, 32'h30000000};
localparam [0:(2**S_WIDTH-1)][31:0]   END_ADDR = {32'h0FFFFFFF, 32'h1FFFFFFF, 32'h2FFFFFFF, 32'h3FFFFFFF};

wire [(2**M_WIDTH-1):0]            M_CLK          ;
wire [(2**M_WIDTH-1):0]            M_RSTN         ;
wire [(2**M_WIDTH-1):0] [M_ID-1:0] M_WR_ADDR_ID   ;
wire [(2**M_WIDTH-1):0] [31:0]     M_WR_ADDR      ;
wire [(2**M_WIDTH-1):0] [ 7:0]     M_WR_ADDR_LEN  ;
wire [(2**M_WIDTH-1):0] [ 1:0]     M_WR_ADDR_BURST;
wire [(2**M_WIDTH-1):0]            M_WR_ADDR_VALID;
wire [(2**M_WIDTH-1):0]            M_WR_ADDR_READY;
wire [(2**M_WIDTH-1):0] [31:0]     M_WR_DATA      ;
wire [(2**M_WIDTH-1):0] [ 3:0]     M_WR_STRB      ;
wire [(2**M_WIDTH-1):0]            M_WR_DATA_LAST ;
wire [(2**M_WIDTH-1):0]            M_WR_DATA_VALID;
wire [(2**M_WIDTH-1):0]            M_WR_DATA_READY;
wire [(2**M_WIDTH-1):0] [M_ID-1:0] M_WR_BACK_ID   ;
wire [(2**M_WIDTH-1):0] [ 1:0]     M_WR_BACK_RESP ;
wire [(2**M_WIDTH-1):0]            M_WR_BACK_VALID;
wire [(2**M_WIDTH-1):0]            M_WR_BACK_READY;
wire [(2**M_WIDTH-1):0] [M_ID-1:0] M_RD_ADDR_ID   ;
wire [(2**M_WIDTH-1):0] [31:0]     M_RD_ADDR      ;
wire [(2**M_WIDTH-1):0] [ 7:0]     M_RD_ADDR_LEN  ;
wire [(2**M_WIDTH-1):0] [ 1:0]     M_RD_ADDR_BURST;
wire [(2**M_WIDTH-1):0]            M_RD_ADDR_VALID;
wire [(2**M_WIDTH-1):0]            M_RD_ADDR_READY;
wire [(2**M_WIDTH-1):0] [M_ID-1:0] M_RD_BACK_ID   ;
wire [(2**M_WIDTH-1):0] [31:0]     M_RD_DATA      ;
wire [(2**M_WIDTH-1):0] [ 1:0]     M_RD_DATA_RESP ;
wire [(2**M_WIDTH-1):0]            M_RD_DATA_LAST ;
wire [(2**M_WIDTH-1):0]            M_RD_DATA_VALID;
wire [(2**M_WIDTH-1):0]            M_RD_DATA_READY;

wire [(2**S_WIDTH-1):0]                    S_CLK          ;
wire [(2**S_WIDTH-1):0]                    S_RSTN         ;
wire [(2**S_WIDTH-1):0] [M_ID+M_WIDTH-1:0] S_WR_ADDR_ID   ;
wire [(2**S_WIDTH-1):0] [31:0]             S_WR_ADDR      ;
wire [(2**S_WIDTH-1):0] [ 7:0]             S_WR_ADDR_LEN  ;
wire [(2**S_WIDTH-1):0] [ 1:0]             S_WR_ADDR_BURST;
wire [(2**S_WIDTH-1):0]                    S_WR_ADDR_VALID;
wire [(2**S_WIDTH-1):0]                    S_WR_ADDR_READY;
wire [(2**S_WIDTH-1):0] [31:0]             S_WR_DATA      ;
wire [(2**S_WIDTH-1):0] [ 3:0]             S_WR_STRB      ;
wire [(2**S_WIDTH-1):0]                    S_WR_DATA_LAST ;
wire [(2**S_WIDTH-1):0]                    S_WR_DATA_VALID;
wire [(2**S_WIDTH-1):0]                    S_WR_DATA_READY;
wire [(2**S_WIDTH-1):0] [M_ID+M_WIDTH-1:0] S_WR_BACK_ID   ;
wire [(2**S_WIDTH-1):0] [ 1:0]             S_WR_BACK_RESP ;
wire [(2**S_WIDTH-1):0]                    S_WR_BACK_VALID;
wire [(2**S_WIDTH-1):0]                    S_WR_BACK_READY;
wire [(2**S_WIDTH-1):0] [M_ID+M_WIDTH-1:0] S_RD_ADDR_ID   ;
wire [(2**S_WIDTH-1):0] [31:0]             S_RD_ADDR      ;
wire [(2**S_WIDTH-1):0] [ 7:0]             S_RD_ADDR_LEN  ;
wire [(2**S_WIDTH-1):0] [ 1:0]             S_RD_ADDR_BURST;
wire [(2**S_WIDTH-1):0]                    S_RD_ADDR_VALID;
wire [(2**S_WIDTH-1):0]                    S_RD_ADDR_READY;
wire [(2**S_WIDTH-1):0] [M_ID+M_WIDTH-1:0] S_RD_BACK_ID   ;
wire [(2**S_WIDTH-1):0] [31:0]             S_RD_DATA      ;
wire [(2**S_WIDTH-1):0] [ 1:0]             S_RD_DATA_RESP ;
wire [(2**S_WIDTH-1):0]                    S_RD_DATA_LAST ;
wire [(2**S_WIDTH-1):0]                    S_RD_DATA_VALID;
wire [(2**S_WIDTH-1):0]                    S_RD_DATA_READY;

wire [0:(2**M_WIDTH-1)] [4:0] M_fifo_empty_flag;
wire [0:(2**S_WIDTH-1)] [4:0] S_fifo_empty_flag;

reg ru_clk;
reg ru_rstn;
// outports wire
wire        	spi_cs;
wire            spi_dq1;
wire        	spi_dq0;
initial ru_clk = 0;
always #50 ru_clk = ~ru_clk;
initial begin
    ru_rstn = 0;
    #10000
    ru_rstn = 1;
end

always #8  BUS_CLK = ~BUS_CLK; //speed:2

initial begin
    BUS_CLK = 0; BUS_RSTN = 0;
#50000
#5000
    BUS_RSTN = 1;
end

integer j;
initial begin
    #5000
    while(~BUS_RSTN) #300;
    while(~S_RSTN[0]) #300;
    #300 M0.set_rd_data_channel(7);
    #300 M0.set_wr_data_channel(1);



    #100000
    #10000 M0.send_rd_addr(2'b00, 32'h00000000, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000001, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000002, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000003, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000004, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000006, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000007, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000008, 8'd000, 2'b00);
    #10000 M0.send_rd_addr(2'b00, 32'h00000009, 8'd000, 2'b00);

    #10000 M0.send_wr_addr(2'b00, 32'h00000000, 8'd000, 2'b00);
    #10000 M0.send_wr_data({16'd10, 1'b1, 3'b000, 12'd123}, 4'b1111);
   
    #1000000
    for(j=0;j<16'd10*4;j=j+1) begin
        #300 M0.send_wr_addr(2'b00, 32'h00000001, 8'd255, 2'b00);
        #300 M0.send_wr_data(j*256, 4'b1111);
    end

    #1000000
    #10000 M0.send_wr_addr(2'b00, 32'h00000004, 8'd000, 2'b00);
    #10000 M0.send_wr_data({31'b0,1'b1}, 4'b1111);
    #10000 M0.send_wr_addr(2'b00, 32'h00000003, 8'd000, 2'b00);
    #10000 M0.send_wr_data({16'd16, 1'b1, 3'b000, 12'd120}, 4'b1111);
    #1000000
    for(j=0;j<16'd16*4;j=j+1) begin
        #300 M0.send_rd_addr(2'b00, 32'h00000005, 8'd255, 2'b00);
    end

end

axi_master_sim M0(
    .MASTER_CLK           (M_CLK [0]        ),
    .MASTER_RSTN          (M_RSTN[0]        ),
    .MASTER_WR_ADDR_ID    (M_WR_ADDR_ID   [0] ),
    .MASTER_WR_ADDR       (M_WR_ADDR      [0] ),
    .MASTER_WR_ADDR_LEN   (M_WR_ADDR_LEN  [0] ),
    .MASTER_WR_ADDR_BURST (M_WR_ADDR_BURST[0] ),
    .MASTER_WR_ADDR_VALID (M_WR_ADDR_VALID[0] ),
    .MASTER_WR_ADDR_READY (M_WR_ADDR_READY[0] ),
    .MASTER_WR_DATA       (M_WR_DATA      [0] ),
    .MASTER_WR_STRB       (M_WR_STRB      [0] ),
    .MASTER_WR_DATA_LAST  (M_WR_DATA_LAST [0] ),
    .MASTER_WR_DATA_VALID (M_WR_DATA_VALID[0] ),
    .MASTER_WR_DATA_READY (M_WR_DATA_READY[0] ),
    .MASTER_WR_BACK_ID    (M_WR_BACK_ID   [0] ),
    .MASTER_WR_BACK_RESP  (M_WR_BACK_RESP [0] ),
    .MASTER_WR_BACK_VALID (M_WR_BACK_VALID[0] ),
    .MASTER_WR_BACK_READY (M_WR_BACK_READY[0] ),
    .MASTER_RD_ADDR_ID    (M_RD_ADDR_ID   [0] ),
    .MASTER_RD_ADDR       (M_RD_ADDR      [0] ),
    .MASTER_RD_ADDR_LEN   (M_RD_ADDR_LEN  [0] ),
    .MASTER_RD_ADDR_BURST (M_RD_ADDR_BURST[0] ),
    .MASTER_RD_ADDR_VALID (M_RD_ADDR_VALID[0] ),
    .MASTER_RD_ADDR_READY (M_RD_ADDR_READY[0] ),
    .MASTER_RD_BACK_ID    (M_RD_BACK_ID   [0] ),
    .MASTER_RD_DATA       (M_RD_DATA      [0] ),
    .MASTER_RD_DATA_RESP  (M_RD_DATA_RESP [0] ),
    .MASTER_RD_DATA_LAST  (M_RD_DATA_LAST [0] ),
    .MASTER_RD_DATA_VALID (M_RD_DATA_VALID[0] ),
    .MASTER_RD_DATA_READY (M_RD_DATA_READY[0] )
);

axi_master_default M1(
    .clk                  (BUS_CLK          ),
    .rstn                 (BUS_RSTN         ),
    .MASTER_CLK           (M_CLK          [1] ),
    .MASTER_RSTN          (M_RSTN         [1] ),
    .MASTER_WR_ADDR_ID    (M_WR_ADDR_ID   [1] ),
    .MASTER_WR_ADDR       (M_WR_ADDR      [1] ),
    .MASTER_WR_ADDR_LEN   (M_WR_ADDR_LEN  [1] ),
    .MASTER_WR_ADDR_BURST (M_WR_ADDR_BURST[1] ),
    .MASTER_WR_ADDR_VALID (M_WR_ADDR_VALID[1] ),
    .MASTER_WR_ADDR_READY (M_WR_ADDR_READY[1] ),
    .MASTER_WR_DATA       (M_WR_DATA      [1] ),
    .MASTER_WR_STRB       (M_WR_STRB      [1] ),
    .MASTER_WR_DATA_LAST  (M_WR_DATA_LAST [1] ),
    .MASTER_WR_DATA_VALID (M_WR_DATA_VALID[1] ),
    .MASTER_WR_DATA_READY (M_WR_DATA_READY[1] ),
    .MASTER_WR_BACK_ID    (M_WR_BACK_ID   [1] ),
    .MASTER_WR_BACK_RESP  (M_WR_BACK_RESP [1] ),
    .MASTER_WR_BACK_VALID (M_WR_BACK_VALID[1] ),
    .MASTER_WR_BACK_READY (M_WR_BACK_READY[1] ),
    .MASTER_RD_ADDR_ID    (M_RD_ADDR_ID   [1] ),
    .MASTER_RD_ADDR       (M_RD_ADDR      [1] ),
    .MASTER_RD_ADDR_LEN   (M_RD_ADDR_LEN  [1] ),
    .MASTER_RD_ADDR_BURST (M_RD_ADDR_BURST[1] ),
    .MASTER_RD_ADDR_VALID (M_RD_ADDR_VALID[1] ),
    .MASTER_RD_ADDR_READY (M_RD_ADDR_READY[1] ),
    .MASTER_RD_BACK_ID    (M_RD_BACK_ID   [1] ),
    .MASTER_RD_DATA       (M_RD_DATA      [1] ),
    .MASTER_RD_DATA_RESP  (M_RD_DATA_RESP [1] ),
    .MASTER_RD_DATA_LAST  (M_RD_DATA_LAST [1] ),
    .MASTER_RD_DATA_VALID (M_RD_DATA_VALID[1] ),
    .MASTER_RD_DATA_READY (M_RD_DATA_READY[1] )
);

axi_master_default M2(
    .clk                  (BUS_CLK           ),
    .rstn                 (BUS_RSTN          ),
    .MASTER_CLK           (M_CLK          [2] ),
    .MASTER_RSTN          (M_RSTN         [2] ),
    .MASTER_WR_ADDR_ID    (M_WR_ADDR_ID   [2] ),
    .MASTER_WR_ADDR       (M_WR_ADDR      [2] ),
    .MASTER_WR_ADDR_LEN   (M_WR_ADDR_LEN  [2] ),
    .MASTER_WR_ADDR_BURST (M_WR_ADDR_BURST[2] ),
    .MASTER_WR_ADDR_VALID (M_WR_ADDR_VALID[2] ),
    .MASTER_WR_ADDR_READY (M_WR_ADDR_READY[2] ),
    .MASTER_WR_DATA       (M_WR_DATA      [2] ),
    .MASTER_WR_STRB       (M_WR_STRB      [2] ),
    .MASTER_WR_DATA_LAST  (M_WR_DATA_LAST [2] ),
    .MASTER_WR_DATA_VALID (M_WR_DATA_VALID[2] ),
    .MASTER_WR_DATA_READY (M_WR_DATA_READY[2] ),
    .MASTER_WR_BACK_ID    (M_WR_BACK_ID   [2] ),
    .MASTER_WR_BACK_RESP  (M_WR_BACK_RESP [2] ),
    .MASTER_WR_BACK_VALID (M_WR_BACK_VALID[2] ),
    .MASTER_WR_BACK_READY (M_WR_BACK_READY[2] ),
    .MASTER_RD_ADDR_ID    (M_RD_ADDR_ID   [2] ),
    .MASTER_RD_ADDR       (M_RD_ADDR      [2] ),
    .MASTER_RD_ADDR_LEN   (M_RD_ADDR_LEN  [2] ),
    .MASTER_RD_ADDR_BURST (M_RD_ADDR_BURST[2] ),
    .MASTER_RD_ADDR_VALID (M_RD_ADDR_VALID[2] ),
    .MASTER_RD_ADDR_READY (M_RD_ADDR_READY[2] ),
    .MASTER_RD_BACK_ID    (M_RD_BACK_ID   [2] ),
    .MASTER_RD_DATA       (M_RD_DATA      [2] ),
    .MASTER_RD_DATA_RESP  (M_RD_DATA_RESP [2] ),
    .MASTER_RD_DATA_LAST  (M_RD_DATA_LAST [2] ),
    .MASTER_RD_DATA_VALID (M_RD_DATA_VALID[2] ),
    .MASTER_RD_DATA_READY (M_RD_DATA_READY[2] )
);

axi_master_default M3(
    .clk                  (BUS_CLK           ),
    .rstn                 (BUS_RSTN          ),
    .MASTER_CLK           (M_CLK          [3] ),
    .MASTER_RSTN          (M_RSTN         [3] ),
    .MASTER_WR_ADDR_ID    (M_WR_ADDR_ID   [3] ),
    .MASTER_WR_ADDR       (M_WR_ADDR      [3] ),
    .MASTER_WR_ADDR_LEN   (M_WR_ADDR_LEN  [3] ),
    .MASTER_WR_ADDR_BURST (M_WR_ADDR_BURST[3] ),
    .MASTER_WR_ADDR_VALID (M_WR_ADDR_VALID[3] ),
    .MASTER_WR_ADDR_READY (M_WR_ADDR_READY[3] ),
    .MASTER_WR_DATA       (M_WR_DATA      [3] ),
    .MASTER_WR_STRB       (M_WR_STRB      [3] ),
    .MASTER_WR_DATA_LAST  (M_WR_DATA_LAST [3] ),
    .MASTER_WR_DATA_VALID (M_WR_DATA_VALID[3] ),
    .MASTER_WR_DATA_READY (M_WR_DATA_READY[3] ),
    .MASTER_WR_BACK_ID    (M_WR_BACK_ID   [3] ),
    .MASTER_WR_BACK_RESP  (M_WR_BACK_RESP [3] ),
    .MASTER_WR_BACK_VALID (M_WR_BACK_VALID[3] ),
    .MASTER_WR_BACK_READY (M_WR_BACK_READY[3] ),
    .MASTER_RD_ADDR_ID    (M_RD_ADDR_ID   [3] ),
    .MASTER_RD_ADDR       (M_RD_ADDR      [3] ),
    .MASTER_RD_ADDR_LEN   (M_RD_ADDR_LEN  [3] ),
    .MASTER_RD_ADDR_BURST (M_RD_ADDR_BURST[3] ),
    .MASTER_RD_ADDR_VALID (M_RD_ADDR_VALID[3] ),
    .MASTER_RD_ADDR_READY (M_RD_ADDR_READY[3] ),
    .MASTER_RD_BACK_ID    (M_RD_BACK_ID   [3] ),
    .MASTER_RD_DATA       (M_RD_DATA      [3] ),
    .MASTER_RD_DATA_RESP  (M_RD_DATA_RESP [3] ),
    .MASTER_RD_DATA_LAST  (M_RD_DATA_LAST [3] ),
    .MASTER_RD_DATA_VALID (M_RD_DATA_VALID[3] ),
    .MASTER_RD_DATA_READY (M_RD_DATA_READY[3] )
);

remote_update_axi_slave #(
    .OFFSET_ADDR            (START_ADDR[0]        ),
	.FPGA_VERSION          	( 48'h2024_1119_1943  ),
	.DEVICE               	( "PG2L100H"          ),
	.USER_BITSTREAM_CNT   	( 2'd3                ),
	.USER_BITSTREAM1_ADDR 	( 24'h40_0000         ),
	.USER_BITSTREAM2_ADDR 	( 24'h80_0000         ),
	.USER_BITSTREAM3_ADDR 	( 24'hC0_0000         ))
S0(
	.clk                 	( ru_clk            ),
	.rstn                	( ru_rstn           ),
	.spi_cs              	( spi_cs            ),
	.spi_dq1             	( spi_dq1           ),
	.spi_dq0             	( spi_dq0           ),
	.SLAVE_CLK           	( S_CLK          [0]  ),
	.SLAVE_RSTN          	( S_RSTN         [0]  ),
	.SLAVE_WR_ADDR_ID    	( S_WR_ADDR_ID   [0]  ),
	.SLAVE_WR_ADDR       	( S_WR_ADDR      [0]  ),
	.SLAVE_WR_ADDR_LEN   	( S_WR_ADDR_LEN  [0]  ),
	.SLAVE_WR_ADDR_BURST 	( S_WR_ADDR_BURST[0]  ),
	.SLAVE_WR_ADDR_VALID 	( S_WR_ADDR_VALID[0]  ),
	.SLAVE_WR_ADDR_READY 	( S_WR_ADDR_READY[0]  ),
	.SLAVE_WR_DATA       	( S_WR_DATA      [0]  ),
	.SLAVE_WR_STRB       	( S_WR_STRB      [0]  ),
	.SLAVE_WR_DATA_LAST  	( S_WR_DATA_LAST [0]  ),
	.SLAVE_WR_DATA_VALID 	( S_WR_DATA_VALID[0]  ),
	.SLAVE_WR_DATA_READY 	( S_WR_DATA_READY[0]  ),
	.SLAVE_WR_BACK_ID    	( S_WR_BACK_ID   [0]  ),
	.SLAVE_WR_BACK_RESP  	( S_WR_BACK_RESP [0]  ),
	.SLAVE_WR_BACK_VALID 	( S_WR_BACK_VALID[0]  ),
	.SLAVE_WR_BACK_READY 	( S_WR_BACK_READY[0]  ),
	.SLAVE_RD_ADDR_ID    	( S_RD_ADDR_ID   [0]  ),
	.SLAVE_RD_ADDR       	( S_RD_ADDR      [0]  ),
	.SLAVE_RD_ADDR_LEN   	( S_RD_ADDR_LEN  [0]  ),
	.SLAVE_RD_ADDR_BURST 	( S_RD_ADDR_BURST[0]  ),
	.SLAVE_RD_ADDR_VALID 	( S_RD_ADDR_VALID[0]  ),
	.SLAVE_RD_ADDR_READY 	( S_RD_ADDR_READY[0]  ),
	.SLAVE_RD_BACK_ID    	( S_RD_BACK_ID   [0]  ),
	.SLAVE_RD_DATA       	( S_RD_DATA      [0]  ),
	.SLAVE_RD_DATA_RESP  	( S_RD_DATA_RESP [0]  ),
	.SLAVE_RD_DATA_LAST  	( S_RD_DATA_LAST [0]  ),
	.SLAVE_RD_DATA_VALID 	( S_RD_DATA_VALID[0]  ),
	.SLAVE_RD_DATA_READY 	( S_RD_DATA_READY[0]  )
);


assign S1_WR_ADDR_READY = 0;assign S2_WR_ADDR_READY = 0;assign S3_WR_ADDR_READY = 0;
assign S1_WR_DATA_READY = 0;assign S2_WR_DATA_READY = 0;assign S3_WR_DATA_READY = 0;
assign S1_WR_BACK_ID    = 0;assign S2_WR_BACK_ID    = 0;assign S3_WR_BACK_ID    = 0;
assign S1_WR_BACK_RESP  = 0;assign S2_WR_BACK_RESP  = 0;assign S3_WR_BACK_RESP  = 0;
assign S1_WR_BACK_VALID = 0;assign S2_WR_BACK_VALID = 0;assign S3_WR_BACK_VALID = 0;
assign S1_RD_ADDR_READY = 0;assign S2_RD_ADDR_READY = 0;assign S3_RD_ADDR_READY = 0;
assign S1_RD_BACK_ID    = 0;assign S2_RD_BACK_ID    = 0;assign S3_RD_BACK_ID    = 0;
assign S1_RD_DATA       = 0;assign S2_RD_DATA       = 0;assign S3_RD_DATA       = 0;
assign S1_RD_DATA_RESP  = 0;assign S2_RD_DATA_RESP  = 0;assign S3_RD_DATA_RESP  = 0;
assign S1_RD_DATA_LAST  = 0;assign S2_RD_DATA_LAST  = 0;assign S3_RD_DATA_LAST  = 0;
assign S1_RD_DATA_VALID = 0;assign S2_RD_DATA_VALID = 0;assign S3_RD_DATA_VALID = 0;

axi_bus #(
	.M_ID       	( M_ID      ),
	.M_WIDTH    	( M_WIDTH   ),
	.S_WIDTH    	( S_WIDTH   ),
	.START_ADDR 	( START_ADDR),
	.END_ADDR   	( END_ADDR  ))
u_axi_bus(
	.BUS_CLK              	( BUS_CLK          ),
	.BUS_RSTN             	( BUS_RSTN         ),
	.MASTER_CLK           	( M_CLK            ),
	.MASTER_RSTN          	( M_RSTN           ),
	.MASTER_WR_ADDR_ID    	( M_WR_ADDR_ID     ),
	.MASTER_WR_ADDR       	( M_WR_ADDR        ),
	.MASTER_WR_ADDR_LEN   	( M_WR_ADDR_LEN    ),
	.MASTER_WR_ADDR_BURST 	( M_WR_ADDR_BURST  ),
	.MASTER_WR_ADDR_VALID 	( M_WR_ADDR_VALID  ),
	.MASTER_WR_ADDR_READY 	( M_WR_ADDR_READY  ),
	.MASTER_WR_DATA       	( M_WR_DATA        ),
	.MASTER_WR_STRB       	( M_WR_STRB        ),
	.MASTER_WR_DATA_LAST  	( M_WR_DATA_LAST   ),
	.MASTER_WR_DATA_VALID 	( M_WR_DATA_VALID  ),
	.MASTER_WR_DATA_READY 	( M_WR_DATA_READY  ),
	.MASTER_WR_BACK_ID    	( M_WR_BACK_ID     ),
	.MASTER_WR_BACK_RESP  	( M_WR_BACK_RESP   ),
	.MASTER_WR_BACK_VALID 	( M_WR_BACK_VALID  ),
	.MASTER_WR_BACK_READY 	( M_WR_BACK_READY  ),
	.MASTER_RD_ADDR_ID    	( M_RD_ADDR_ID     ),
	.MASTER_RD_ADDR       	( M_RD_ADDR        ),
	.MASTER_RD_ADDR_LEN   	( M_RD_ADDR_LEN    ),
	.MASTER_RD_ADDR_BURST 	( M_RD_ADDR_BURST  ),
	.MASTER_RD_ADDR_VALID 	( M_RD_ADDR_VALID  ),
	.MASTER_RD_ADDR_READY 	( M_RD_ADDR_READY  ),
	.MASTER_RD_BACK_ID    	( M_RD_BACK_ID     ),
	.MASTER_RD_DATA       	( M_RD_DATA        ),
	.MASTER_RD_DATA_RESP  	( M_RD_DATA_RESP   ),
	.MASTER_RD_DATA_LAST  	( M_RD_DATA_LAST   ),
	.MASTER_RD_DATA_VALID 	( M_RD_DATA_VALID  ),
	.MASTER_RD_DATA_READY 	( M_RD_DATA_READY  ),
	.SLAVE_CLK            	( S_CLK            ),
	.SLAVE_RSTN           	( S_RSTN           ),
	.SLAVE_WR_ADDR_ID     	( S_WR_ADDR_ID     ),
	.SLAVE_WR_ADDR        	( S_WR_ADDR        ),
	.SLAVE_WR_ADDR_LEN    	( S_WR_ADDR_LEN    ),
	.SLAVE_WR_ADDR_BURST  	( S_WR_ADDR_BURST  ),
	.SLAVE_WR_ADDR_VALID  	( S_WR_ADDR_VALID  ),
	.SLAVE_WR_ADDR_READY  	( S_WR_ADDR_READY  ),
	.SLAVE_WR_DATA        	( S_WR_DATA        ),
	.SLAVE_WR_STRB        	( S_WR_STRB        ),
	.SLAVE_WR_DATA_LAST   	( S_WR_DATA_LAST   ),
	.SLAVE_WR_DATA_VALID  	( S_WR_DATA_VALID  ),
	.SLAVE_WR_DATA_READY  	( S_WR_DATA_READY  ),
	.SLAVE_WR_BACK_ID     	( S_WR_BACK_ID     ),
	.SLAVE_WR_BACK_RESP   	( S_WR_BACK_RESP   ),
	.SLAVE_WR_BACK_VALID  	( S_WR_BACK_VALID  ),
	.SLAVE_WR_BACK_READY  	( S_WR_BACK_READY  ),
	.SLAVE_RD_ADDR_ID     	( S_RD_ADDR_ID     ),
	.SLAVE_RD_ADDR        	( S_RD_ADDR        ),
	.SLAVE_RD_ADDR_LEN    	( S_RD_ADDR_LEN    ),
	.SLAVE_RD_ADDR_BURST  	( S_RD_ADDR_BURST  ),
	.SLAVE_RD_ADDR_VALID  	( S_RD_ADDR_VALID  ),
	.SLAVE_RD_ADDR_READY  	( S_RD_ADDR_READY  ),
	.SLAVE_RD_BACK_ID     	( S_RD_BACK_ID     ),
	.SLAVE_RD_DATA        	( S_RD_DATA        ),
	.SLAVE_RD_DATA_RESP   	( S_RD_DATA_RESP   ),
	.SLAVE_RD_DATA_LAST   	( S_RD_DATA_LAST   ),
	.SLAVE_RD_DATA_VALID  	( S_RD_DATA_VALID  ),
	.SLAVE_RD_DATA_READY  	( S_RD_DATA_READY  ),
	.M_fifo_empty_flag    	( M_fifo_empty_flag),
	.S_fifo_empty_flag    	( S_fifo_empty_flag)
);

reg grs_n;
GTP_GRS GRS_INST(.GRS_N (grs_n));
initial begin
grs_n = 1'b0;
#5 grs_n = 1'b1;
end

MX25L12805D flash_u( ru_clk, spi_cs, spi_dq0, spi_dq1, 1'b0, 1'b1 );


endmodule