module led_display_in_axi_slave (
    input clk,
    input rstn,
    input sck,
    input ser,
    input rck,

    output wire         SLAVE_CLK          ,
    output wire         SLAVE_RSTN         ,

    input  wire [4-1:0] SLAVE_WR_ADDR_ID   ,
    input  wire [31:0]  SLAVE_WR_ADDR      ,
    input  wire [ 7:0]  SLAVE_WR_ADDR_LEN  ,
    input  wire [ 1:0]  SLAVE_WR_ADDR_BURST,
    input  wire         SLAVE_WR_ADDR_VALID,
    output wire         SLAVE_WR_ADDR_READY,

    input  wire [31:0]  SLAVE_WR_DATA      ,
    input  wire [ 3:0]  SLAVE_WR_STRB      ,
    input  wire         SLAVE_WR_DATA_LAST ,
    input  wire         SLAVE_WR_DATA_VALID,
    output wire         SLAVE_WR_DATA_READY,

    output wire [4-1:0] SLAVE_WR_BACK_ID   ,
    output wire [ 1:0]  SLAVE_WR_BACK_RESP ,
    output wire         SLAVE_WR_BACK_VALID,
    input  wire         SLAVE_WR_BACK_READY,

    input  wire [4-1:0] SLAVE_RD_ADDR_ID   ,
    input  wire [31:0]  SLAVE_RD_ADDR      ,
    input  wire [ 7:0]  SLAVE_RD_ADDR_LEN  ,
    input  wire [ 1:0]  SLAVE_RD_ADDR_BURST,
    input  wire         SLAVE_RD_ADDR_VALID,
    output wire         SLAVE_RD_ADDR_READY,
    output wire [4-1:0] SLAVE_RD_BACK_ID   ,

    output wire [31:0]  SLAVE_RD_DATA      ,
    output wire [ 1:0]  SLAVE_RD_DATA_RESP ,
    output wire         SLAVE_RD_DATA_LAST ,
    output wire         SLAVE_RD_DATA_VALID,
    input  wire         SLAVE_RD_DATA_READY
);
//只能读
rstn_sync led_display_rstn_sync(clk,rstn,SLAVE_RSTN);
assign SLAVE_CLK = clk;
assign SLAVE_WR_ADDR_READY = 0;
assign SLAVE_WR_DATA_READY = 0;
assign SLAVE_WR_BACK_ID    = 0;
assign SLAVE_WR_BACK_RESP  = 0;
assign SLAVE_WR_BACK_VALID = 0;
//****************************************************//
wire QS;
wire [7:0] led_display_in_seg;
wire [31:0] led_display_in_sel;
wire [4:0] decoder_in;//5bit
SIM_74HC595  SIM_74HC595_inst_seg (
    .sck(sck),
    .rstn(SLAVE_RSTN),
    .rck(rck),
    .ser(ser),
    .QS(QS),
    .out(led_display_in_seg)
  );
SIM_74HC595  SIM_74HC595_inst_sel (
    .sck(sck),
    .rstn(SLAVE_RSTN),
    .rck(rck),
    .ser(QS),
    .QS(),
    .out(decoder_in)
  );
decoder_5_32  decoder_5_32_inst (
    .in(decoder_in),
    .sel(led_display_in_sel)
  );
reg [7:0] led [31:0];
integer i;
always @(posedge clk or negedge SLAVE_RSTN) begin
    if (~SLAVE_RSTN) begin
        for (i = 0; i < 32; i = i + 1) 
            led[i] <= 8'd0;
    end else begin
        for (i = 0; i < 32; i = i + 1) begin
            if (led_display_in_sel[i]) 
                led[i] <= led_display_in_seg;
        end
    end
end
//****************************************************//
reg rd_en;
reg [ 7:0] txcnt    ;
reg [ 3:0] rdaddrid ;
reg [31:0] rdaddr   ;
reg [ 7:0] rdaddrlen;
reg [31:0] rddata   ;
assign SLAVE_RD_BACK_ID = rdaddrid;
assign SLAVE_RD_ADDR_READY = ~rd_en;
always @(posedge clk or SLAVE_RSTN) begin
    if(~SLAVE_RSTN)begin
        rdaddrid  <= 'd0;
        rdaddrlen <= 'd0;
    end
    else if(SLAVE_RD_ADDR_VALID && SLAVE_RD_ADDR_READY)begin
        rdaddrid  <= SLAVE_RD_ADDR_ID;
        rdaddrlen <= SLAVE_RD_ADDR_LEN;
    end
    else begin
        rdaddrid  <= rdaddrid ;
        rdaddrlen <= rdaddrlen;
    end
end
always @(posedge clk or negedge SLAVE_RSTN) begin
    if(~SLAVE_RSTN) rdaddr <= 'd0;
    else if(SLAVE_RD_ADDR_VALID && SLAVE_RD_ADDR_READY) rdaddr <= SLAVE_RD_ADDR;
    else if(SLAVE_RD_DATA_VALID && SLAVE_RD_DATA_READY && ~SLAVE_RD_DATA_LAST) rdaddr <= rdaddr + 1;
    else rdaddr <= rdaddr;
end
always @(posedge clk or negedge SLAVE_RSTN) begin
    if(~SLAVE_RSTN) rd_en <= 0;
    else if(SLAVE_RD_ADDR_VALID && SLAVE_RD_ADDR_READY) rd_en <= 1;
    else if(SLAVE_RD_DATA_VALID && SLAVE_RD_DATA_READY && SLAVE_RD_DATA_LAST) rd_en <= 0;
    else rd_en <= rd_en;
end
always @(posedge clk or negedge SLAVE_RSTN) begin
    if(~SLAVE_RSTN) txcnt <= 0;
    else if(SLAVE_RD_ADDR_VALID && SLAVE_RD_ADDR_READY) txcnt <= 0;
    else if(SLAVE_RD_DATA_VALID && SLAVE_RD_DATA_READY) begin
        if(~SLAVE_RD_DATA_LAST)
            txcnt <= txcnt + 1;
        else 
            txcnt <= 0;
    end
    else txcnt <= txcnt;
end
assign SLAVE_RD_DATA_VALID = rd_en;
assign SLAVE_RD_DATA       = rddata;
assign SLAVE_RD_DATA_RESP  = rddata < 32'd32 ? 2'b00 : 2'b10;
assign SLAVE_RD_DATA_LAST  = txcnt == rdaddrlen ? 1'b1 : 1'b0;
always @(*) begin
    case(rdaddr)
        32'd0  : rddata = {19'd0 , 5'd0  , led[0 ]};
        32'd1  : rddata = {19'd0 , 5'd1  , led[1 ]};
        32'd2  : rddata = {19'd0 , 5'd2  , led[2 ]};
        32'd3  : rddata = {19'd0 , 5'd3  , led[3 ]};
        32'd4  : rddata = {19'd0 , 5'd4  , led[4 ]};
        32'd5  : rddata = {19'd0 , 5'd5  , led[5 ]};
        32'd6  : rddata = {19'd0 , 5'd6  , led[6 ]};
        32'd7  : rddata = {19'd0 , 5'd7  , led[7 ]};
        32'd8  : rddata = {19'd0 , 5'd8  , led[8 ]};
        32'd9  : rddata = {19'd0 , 5'd9  , led[9 ]};
        32'd10 : rddata = {19'd0 , 5'd10 , led[10]};
        32'd11 : rddata = {19'd0 , 5'd11 , led[11]};
        32'd12 : rddata = {19'd0 , 5'd12 , led[12]};
        32'd13 : rddata = {19'd0 , 5'd13 , led[13]};
        32'd14 : rddata = {19'd0 , 5'd14 , led[14]};
        32'd15 : rddata = {19'd0 , 5'd15 , led[15]};
        32'd16 : rddata = {19'd0 , 5'd16 , led[16]};
        32'd17 : rddata = {19'd0 , 5'd17 , led[17]};
        32'd18 : rddata = {19'd0 , 5'd18 , led[18]};
        32'd19 : rddata = {19'd0 , 5'd19 , led[19]};
        32'd20 : rddata = {19'd0 , 5'd20 , led[20]};
        32'd21 : rddata = {19'd0 , 5'd21 , led[21]};
        32'd22 : rddata = {19'd0 , 5'd22 , led[22]};
        32'd23 : rddata = {19'd0 , 5'd23 , led[23]};
        32'd24 : rddata = {19'd0 , 5'd24 , led[24]};
        32'd25 : rddata = {19'd0 , 5'd25 , led[25]};
        32'd26 : rddata = {19'd0 , 5'd26 , led[26]};
        32'd27 : rddata = {19'd0 , 5'd27 , led[27]};
        32'd28 : rddata = {19'd0 , 5'd28 , led[28]};
        32'd29 : rddata = {19'd0 , 5'd29 , led[29]};
        32'd30 : rddata = {19'd0 , 5'd30 , led[30]};
        32'd31 : rddata = {19'd0 , 5'd31 , led[31]};
        default : rddata = 32'hFFFFFFFF;
    endcase
end

endmodule