`timescale  1ns/1ns
////////////////////////////////////////////////////////////////////////
// Author  : EmbedFire
// ʵ��ƽ̨: Ұ��FPGAϵ�п�����
// ��˾    : http://www.embedfire.com
// ��̳    : http://www.firebbs.cn
// �Ա�    : https://fire-stm32.taobao.com
////////////////////////////////////////////////////////////////////////

module udp_tx (
    input                clk        , //ʱ���ź�
    input                rst_n      , //��λ�źţ��͵�ƽ��Ч

    input                tx_start_en/* synthesis PAP_MARK_DEBUG=��true�� */, //��̫����ʼ�����ź�
    input        [31:0]  tx_data    /* synthesis PAP_MARK_DEBUG=��true�� */, //��̫������������
    input        [15:0]  tx_byte_num/* synthesis PAP_MARK_DEBUG=��true�� */, //��̫�����͵���Ч�ֽ���
    input        [31:0]  crc_data   , //CRCУ������
    input         [7:0]  crc_next   , //CRC�´�У���������
    input                udp_tx_sel /* synthesis PAP_MARK_DEBUG=��true�� */,
    output  reg          udp_tx_req /* synthesis PAP_MARK_DEBUG=��true�� */,
    output  reg          udp_tx_working,
    output  reg          tx_done    /* synthesis PAP_MARK_DEBUG=��true�� */, //��̫����������ź�
    output  reg          tx_req     /* synthesis PAP_MARK_DEBUG=��true�� */, //�����������ź�
    output  reg          gmii_tx_en /* synthesis PAP_MARK_DEBUG=��true�� */, //GMII���������Ч�ź�
    output  reg  [7:0]   gmii_txd   /* synthesis PAP_MARK_DEBUG=��true�� */, //GMII�������
    output  reg          crc_en     , //CRC��ʼУ��ʹ��
    output  reg          crc_clr    , //CRC���ݸ�λ�ź�
    input                timestamp_rst,
    input        [31:0]  des_ip   ,
    input        [47:0]  des_mac  ,
    input        [31:0]  board_ip ,
    input        [47:0]  board_mac
    );

localparam  st_wait      = 7'b000_0000; //�ȴ��ٲ�����Ӧ
localparam  st_idle      = 7'b000_0001; //��ʼ״̬���ȴ���ʼ�����ź�
localparam  st_check_sum = 7'b000_0010; //IP�ײ�У���
localparam  st_preamble  = 7'b000_0100; //����ǰ����+֡��ʼ�綨��
localparam  st_eth_head  = 7'b000_1000; //������̫��֡ͷ
localparam  st_ip_head   = 7'b001_0000; //����IP�ײ�+UDP�ײ�
localparam  st_tx_data   = 7'b010_0000; //��������
localparam  st_crc       = 7'b100_0000; //����CRCУ��ֵ

localparam  ETH_TYPE      = 16'h0800  ;  //��̫��Э������ IPЭ��
localparam  SOURCE_PORT   = 16'd1234; //Դ�˿ں�
localparam  DEST_PORT_MIN = 16'd1234; //Ŀ�Ķ˿ںŷ�Χ��Сֵ
localparam  DEST_PORT_MAX = 16'd1244; //Ŀ�Ķ˿ںŷ�Χ���ֵ
//��̫��������С46���ֽڣ�IP�ײ�20���ֽ�+UDP�ײ�8���ֽ�
//������������46-20-8=18���ֽ�
localparam  MIN_DATA_NUM = 16'd18 - 16'd4    ; //����ʱ���4�ֽ�

//reg define
reg  [6:0]   cur_state      /* synthesis PAP_MARK_DEBUG=��true�� */;
reg  [6:0]   next_state     ;

reg  [7:0]   preamble[7:0]  ; //ǰ����
reg  [7:0]   eth_head[13:0] ; //��̫���ײ�
reg  [31:0]  ip_head[7:0]   ; //IP�ײ� + UDP�ײ� + ʱ���(����ip_head[7]����32λʱ���)

reg          start_en_d0    ;
reg          start_en_d1    ;
reg  [15:0]  tx_data_num    ; //���͵���Ч�����ֽڸ���
reg  [15:0]  total_num      ; //���ֽ���
reg          trig_tx_en     ;
reg  [15:0]  udp_num        ; //UDP�ֽ���
reg          skip_en        /* synthesis PAP_MARK_DEBUG=��true�� */; //����״̬��תʹ���ź�
reg  [4:0]   cnt            ;
reg  [31:0]  check_buffer   ; //�ײ�У���
reg  [1:0]   tx_bit_sel     ;
reg  [15:0]  data_cnt       ; //�������ݸ���������
reg          tx_done_t      ;
reg  [4:0]   real_add_cnt   ; //��̫������ʵ�ʶ෢���ֽ���
reg  [15:0]  des_port       ; //Ŀ�Ķ˿ں�
reg  [31:0]  dec_ip_reg     ;

// 32λ��������������ʱ���
reg  [31:0]  packet_counter /* synthesis PAP_MARK_DEBUG="true" */;
//wire define
wire         pos_start_en    ;//��ʼ��������������
wire [15:0]  real_tx_data_num;//ʵ�ʷ��͵��ֽ���(��̫�������ֽ�Ҫ��)
//*****************************************************
//**                    main code
//*****************************************************

always @(*) begin
    eth_head[0]  <= des_mac[47:40];
    eth_head[1]  <= des_mac[39:32];
    eth_head[2]  <= des_mac[31:24];
    eth_head[3]  <= des_mac[23:16];
    eth_head[4]  <= des_mac[15:8];
    eth_head[5]  <= des_mac[7:0];
    eth_head[6]  <= board_mac[47:40];
    eth_head[7]  <= board_mac[39:32];
    eth_head[8]  <= board_mac[31:24];
    eth_head[9]  <= board_mac[23:16];
    eth_head[10] <= board_mac[15:8];
    eth_head[11] <= board_mac[7:0];
    dec_ip_reg   <= des_ip;
end
assign  pos_start_en = (~start_en_d1) & start_en_d0;
assign  real_tx_data_num = ((tx_data_num) >= MIN_DATA_NUM)
                           ? (tx_data_num) : MIN_DATA_NUM;

//��tx_start_en��������
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        start_en_d0 <= 1'b0;
        start_en_d1 <= 1'b0;
    end
    else begin
        start_en_d0 <= tx_start_en;
        start_en_d1 <= start_en_d0;
    end
end

//�Ĵ�������Ч�ֽ�
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        tx_data_num <= 16'd0;
        total_num <= 16'd0;
        udp_num <= 16'd0;
    end
    else begin
        if(pos_start_en && cur_state==st_idle) begin
            //���ݳ��ȣ��������ݣ�
            tx_data_num <= tx_byte_num; //����ʱ���4�ֽ�
            //IP���ȣ���Ч����+IP�ײ�����(20�ֽ�)+UDP�ײ�����(8�ֽ�)
            total_num <= (tx_byte_num + 16'd4) + 16'd28;
            //UDP���ȣ���Ч����+UDP�ײ�����(8�ֽ�)
            udp_num <= (tx_byte_num + 16'd4) + 16'd8;
        end
    end
end

//���������ź�
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        trig_tx_en <= 1'b0;
    else
        trig_tx_en <= pos_start_en;

end

always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cur_state <= st_idle;
    else
        cur_state <= next_state;
end

always @(*) begin
    next_state = st_idle;
    case(cur_state)
        st_idle     : begin                               //�ȴ���������
            if(skip_en)
                next_state = st_wait;
            else
                next_state = st_idle;
        end
        st_wait : begin                                  //�ȴ��ٲ�����Ӧ
            if(skip_en)
                next_state = st_check_sum;
            else
                next_state = st_wait;

        end
        st_check_sum: begin                               //IP�ײ�У��
            if(skip_en)
                next_state = st_preamble;
            else
                next_state = st_check_sum;
        end
        st_preamble : begin                               //����ǰ����+֡��ʼ�綨��
            if(skip_en)
                next_state = st_eth_head;
            else
                next_state = st_preamble;
        end
        st_eth_head : begin                               //������̫���ײ�
            if(skip_en)
                next_state = st_ip_head;
            else
                next_state = st_eth_head;
        end
        st_ip_head : begin                                //����IP�ײ�+UDP�ײ�
            if(skip_en)
                next_state = st_tx_data;
            else
                next_state = st_ip_head;
        end
        st_tx_data : begin                                //��������
            if(skip_en)
                next_state = st_crc;
            else
                next_state = st_tx_data;
        end
        st_crc: begin                                     //����CRCУ��ֵ
            if(skip_en)
                next_state = st_idle;
            else
                next_state = st_crc;
        end
        default : next_state = st_idle;
    endcase
end

//��������
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        skip_en         <= 1'b0;
        cnt             <= 5'd0;
        check_buffer    <= 32'd0;
        ip_head[1][31:16] <= 16'd0;
        tx_bit_sel      <= 2'b0;
        crc_en          <= 1'b0;
        gmii_tx_en      <= 1'b0;
        gmii_txd        <= 8'd0;
        tx_req          <= 1'b0;
        tx_done_t       <= 1'b0;
        data_cnt        <= 16'd0;
        real_add_cnt    <= 5'd0;
        udp_tx_working  <= 0;
        udp_tx_req      <= 0;
        des_port        <= DEST_PORT_MIN; //��ʼ��Ŀ�Ķ˿ں�
        //��ʼ������
        //ǰ���� 7��8'h55 + 1��8'hd5
        preamble[0] <= 8'h55;
        preamble[1] <= 8'h55;
        preamble[2] <= 8'h55;
        preamble[3] <= 8'h55;
        preamble[4] <= 8'h55;
        preamble[5] <= 8'h55;
        preamble[6] <= 8'h55;
        preamble[7] <= 8'hd5;
        //��̫������
        eth_head[12] <= ETH_TYPE[15:8];
        eth_head[13] <= ETH_TYPE[7:0];
    end
    else begin
        skip_en <= 1'b0;
        tx_req <= 1'b0;
        crc_en <= 1'b0;
        gmii_tx_en <= 1'b0;
        tx_done_t <= 1'b0;
        case(next_state)
            st_idle     : begin
                udp_tx_working <= 0;
                if(trig_tx_en) begin
                    skip_en <= 1'b1;
                    //�汾�ţ�4 �ײ����ȣ�5(��λ:32bit,20byte/4=5)
                    ip_head[0] <= {8'h45,8'h00,total_num};
                    //16λ��ʶ��ÿ�η����ۼ�1
                    ip_head[1][31:16] <= ip_head[1][31:16] + 1'b1;
                    //bit[15:13]: 010��ʾ����Ƭ
                    ip_head[1][15:0] <= 16'h4000;
                    //Э�飺17(udp)
                    ip_head[2] <= {8'h40,8'd17,16'h0};
                    //ԴIP��ַ
                    ip_head[3] <= board_ip;
                    //Ŀ��IP��ַ
                    ip_head[4] <= dec_ip_reg;
                    //16λԴ�˿ںţ�1234  16λĿ�Ķ˿ںţ�1234
                    ip_head[5] <= {SOURCE_PORT,des_port};
                    des_port <= (des_port < DEST_PORT_MAX) ? (des_port + 1'b1) : (DEST_PORT_MIN);
                    // des_port <= DEST_PORT_MIN;
                    //16λudp���ȣ�16λudpУ���
                    ip_head[6] <= {udp_num,16'h0000};
                    //32λʱ���
                    ip_head[7] <= packet_counter;
                end
            end
            st_wait : begin
                if(udp_tx_sel)begin
                    udp_tx_working <= 1;
                    skip_en <= 1;
                    udp_tx_req <= 0;
                end
                else begin
                    udp_tx_working <= 0;
                    skip_en <= 0;
                    udp_tx_req <= 1;
                end
            end
            st_check_sum: begin                           //IP�ײ�У��
                cnt <= cnt + 5'd1;
                if(cnt == 5'd0) begin
                    check_buffer <= ip_head[0][31:16] + ip_head[0][15:0]
                                  + ip_head[1][31:16] + ip_head[1][15:0]
                                  + ip_head[2][31:16] + ip_head[2][15:0]
                                  + ip_head[3][31:16] + ip_head[3][15:0]
                                  + ip_head[4][31:16] + ip_head[4][15:0];
                end
                else if(cnt == 5'd1)                      //���ܳ��ֽ�λ,�ۼ�һ��
                    check_buffer <= check_buffer[31:16] + check_buffer[15:0];
                else if(cnt == 5'd2) begin                //�����ٴγ��ֽ�λ,�ۼ�һ��
                    check_buffer <= check_buffer[31:16] + check_buffer[15:0];
                end
                else if(cnt == 5'd3) begin                //��λȡ��
                    skip_en <= 1'b1;
                    cnt <= 5'd0;
                    ip_head[2][15:0] <= ~check_buffer[15:0];
                end
            end
            st_preamble : begin                           //����ǰ����+֡��ʼ�綨��
                gmii_tx_en <= 1'b1;
                gmii_txd <= preamble[cnt];
                if(cnt == 5'd7) begin
                    skip_en <= 1'b1;
                    cnt <= 5'd0;
                end
                else
                    cnt <= cnt + 5'd1;
            end
            st_eth_head : begin                           //������̫���ײ�
                gmii_tx_en <= 1'b1;
                crc_en <= 1'b1;
                gmii_txd <= eth_head[cnt];
                if (cnt == 5'd13) begin
                    skip_en <= 1'b1;
                    cnt <= 5'd0;
                end
                else
                    cnt <= cnt + 5'd1;
            end
            st_ip_head  : begin                           //����IP�ײ� + UDP�ײ� + ʱ���
                crc_en <= 1'b1;
                gmii_tx_en <= 1'b1;
                tx_bit_sel <= tx_bit_sel + 2'd1;
                if(tx_bit_sel == 3'd0)
                    gmii_txd <= ip_head[cnt][31:24];
                else if(tx_bit_sel == 3'd1)
                    gmii_txd <= ip_head[cnt][23:16];
                else if(tx_bit_sel == 3'd2) begin
                    gmii_txd <= ip_head[cnt][15:8];
                    if(cnt == 5'd7) begin
                        //��ǰ���������ݣ��ȴ�������Чʱ����
                        tx_req <= 1'b1;
                    end
                end
                else if(tx_bit_sel == 3'd3) begin
                    gmii_txd <= ip_head[cnt][7:0];
                    if(cnt == 5'd7) begin
                        skip_en <= 1'b1;
                        cnt <= 5'd0;
                    end
                    else
                        cnt <= cnt + 5'd1;
                end
            end
            st_tx_data  : begin                           //��������
                crc_en <= 1'b1;
                gmii_tx_en <= 1'b1;
                tx_bit_sel <= tx_bit_sel + 3'd1;
                if(data_cnt < tx_data_num - 16'd1)
                    data_cnt <= data_cnt + 16'd1;
                else if(data_cnt == tx_data_num - 16'd1)begin
                    //������͵���Ч��������18���ֽڣ��ں������λ
                    //�����ֵΪ���һ�η��͵���Ч����
                    gmii_txd <= 8'd0;
                    if(data_cnt + real_add_cnt < real_tx_data_num - 16'd1)
                        real_add_cnt <= real_add_cnt + 5'd1;
                    else begin
                        skip_en <= 1'b1;
                        data_cnt <= 16'd0;
                        real_add_cnt <= 5'd0;
                        tx_bit_sel <= 3'd0;
                    end
                end
                if(tx_bit_sel == 1'b0)
                    gmii_txd <= tx_data[31:24];
                else if(tx_bit_sel == 3'd1)
                    gmii_txd <= tx_data[23:16];
                else if(tx_bit_sel == 3'd2) begin
                    gmii_txd <= tx_data[15:8];
                    if(data_cnt != tx_data_num - 16'd1 && data_cnt != tx_data_num - 16'd2)
                        tx_req <= 1'b1;
                end
                else if(tx_bit_sel == 3'd3)
                    gmii_txd <= tx_data[7:0];
            end
            st_crc      : begin                          //����CRCУ��ֵ
                gmii_tx_en <= 1'b1;
                tx_bit_sel <= tx_bit_sel + 3'd1;
                if(tx_bit_sel == 3'd0)
                    gmii_txd <= {~crc_next[0], ~crc_next[1], ~crc_next[2],~crc_next[3],
                                 ~crc_next[4], ~crc_next[5], ~crc_next[6],~crc_next[7]};
                else if(tx_bit_sel == 3'd1)
                    gmii_txd <= {~crc_data[16], ~crc_data[17], ~crc_data[18],~crc_data[19],
                                 ~crc_data[20], ~crc_data[21], ~crc_data[22],~crc_data[23]};
                else if(tx_bit_sel == 3'd2) begin
                    gmii_txd <= {~crc_data[8], ~crc_data[9], ~crc_data[10],~crc_data[11],
                                 ~crc_data[12], ~crc_data[13], ~crc_data[14],~crc_data[15]};
                end
                else if(tx_bit_sel == 3'd3) begin
                    gmii_txd <= {~crc_data[0], ~crc_data[1], ~crc_data[2],~crc_data[3],
                                 ~crc_data[4], ~crc_data[5], ~crc_data[6],~crc_data[7]};
                    tx_done_t <= 1'b1;
                    skip_en <= 1'b1;
                end
            end
            default :;
        endcase
    end
end

//��������źż�crcֵ��λ�ź�
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        tx_done <= 1'b0;
        crc_clr <= 1'b0;
    end
    else begin
        tx_done <= tx_done_t;
        crc_clr <= tx_done_t;
    end
end

always @(posedge clk or negedge rst_n) begin
    if(!rst_n) packet_counter <= 32'd0;
    else if(timestamp_rst) packet_counter <= 32'd0;
    else if(tx_done_t) packet_counter <= packet_counter + 1'b1;
    else packet_counter <= packet_counter;
end

endmodule

