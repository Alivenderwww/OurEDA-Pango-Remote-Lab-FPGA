module dso_top #(
    parameter CLK_FS = 32'd50_000_000 // 基准时钟频率值
)(
    input         clk,
    input         rstn,       // 复位信号

    input         ad_clk,     // AD时钟
    input  [7:0]  ad_data,    // AD输入数据

    input         wave_run,   // 波形采集启动/停止
    input  [7:0]  trig_level, // 触发电平
    input         trig_edge,  // 触发边沿
    input  [9:0]  deci_rate,  // 抽样率

    input         ram_refresh/* synthesis PAP_MARK_DEBUG="true" */,
    input  [9:0]  wave_rd_addr/* synthesis PAP_MARK_DEBUG="true" */, // RAM读地址 0-299
    output [7:0]  wave_rd_data/* synthesis PAP_MARK_DEBUG="true" */, // RAM读数据
	output        wave_ready/* synthesis PAP_MARK_DEBUG="true" */,   // RAM读数据准备好
	output [9:0]  wave_trig_addr/* synthesis PAP_MARK_DEBUG="true" */, // 触发地址

    output        outrange,     //水平偏移超出范围
    output        ad_pulse,     //AD采样脉冲
    output [19:0] ad_freq/* synthesis PAP_MARK_DEBUG="true" */,      //AD采样频率
    output [7:0]  ad_vpp/* synthesis PAP_MARK_DEBUG="true" */,       //AD采样幅度
    output [7:0]  ad_max/* synthesis PAP_MARK_DEBUG="true" */,       //AD采样最大值
    output [7:0]  ad_min/* synthesis PAP_MARK_DEBUG="true" */        //AD采样最小值
);

wire       	deci_valid;

//参数测量模块
param_measure #(
	.CLK_FS 	( CLK_FS  ))
u_param_measure(
	.clk        	( clk         ),
	.rstn       	( rstn        ),
	.trig_level 	( trig_level  ),
	.ad_clk     	( ad_clk      ),
	.ad_data    	( ad_data     ),
	.ad_pulse   	( ad_pulse    ),
	.ad_freq    	( ad_freq     ),
	.ad_vpp     	( ad_vpp      ),
	.ad_max     	( ad_max      ),
	.ad_min     	( ad_min      )
);

//数据存储模块
data_store u_data_store(
	.rstn         	( rstn           ),
	.trig_level    	( trig_level     ),
	.trig_edge     	( trig_edge      ),
	.wave_run      	( wave_run       ),
	.ad_clk        	( ad_clk         ),
	.ad_data       	( ad_data        ),
	.deci_valid    	( deci_valid     ),
	.ram_rd_clk     ( clk            ),
	.ram_refresh   	( ram_refresh    ),
	.wave_rd_addr  	( wave_rd_addr   ),
	.wave_rd_data  	( wave_rd_data   ),
    .wave_ready		( wave_ready	 ),
    .wave_trig_addr	( wave_trig_addr )
);

//抽样模块
decimator u_decimator(
	.ad_clk     	( ad_clk      ),
	.rstn       	( rstn        ),
	.deci_rate  	( deci_rate   ),
	.deci_valid 	( deci_valid  )
);


endmodule //dso_top
