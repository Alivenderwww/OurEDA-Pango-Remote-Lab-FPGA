module ws2812_ctrl(

);


endmodule