module data_ctrl_slave #(
parameter OFFSET_ADDR           = 32'h3000_0000     ,
parameter FPGA_VERSION          = 48'h2000_0101_1200    // year,month,day,hour,minute;
)(
input  wire        clk                     ,
input  wire        rstn                    ,

//写入比特流-控制接口
output reg          flash_wr_en             ,
output reg  [11:0]  start_wr_sector     ,
output reg  [15:0]  wr_sector_num           ,
input               flash_wr_done           ,
input               flash_clear_done        ,
//写入比特流-数据接口
output wire        bitstream_fifo_rd_rdy   ,
input  wire        bitstream_fifo_rd_req   ,
output wire        bitstream_valid         ,
output wire [7:0]  bitstream_data          ,
output wire        bitstream_eop           ,

//读出比特流-控制接口1
output reg          flash_rd_en             ,
output reg  [11:0]  start_rd_sub_sector     ,
output reg  [15:0]  rd_sector_num           ,
input               flash_rd_done           ,
//读出比特流-控制接口2
input  wire        bs_readback_crc_valid   ,
input  wire [31:0] bs_readback_crc         ,
//读出比特流-控制接口3
output  reg        crc_check_en            ,
output  reg [1:0]  bs_crc32_ok             ,//[1]:valid   [0]:1'b0,OK  1'b1,error
//读出比特流-回读接口
output  reg        bitstream_up2cpu_en     ,
output wire        flash_rd_data_fifo_afull,
input  wire [7:0]  flash_rd_data           ,
input  wire        flash_rd_valid          ,

//热启动接口
output  reg        hotreset_en             ,
output  reg [23:0] hotreset_addr           ,
//未知用途
input  wire        ipal_busy               ,
input  wire        time_out_reg            ,
//弃用
input  wire [15:0] flash_flag_status       ,
output wire        flash_cfg_cmd_en        ,
output wire [7:0]  flash_cfg_cmd           ,
output wire [15:0] flash_cfg_reg_wrdata    ,
input  wire        flash_cfg_reg_rd_en     ,
input  wire [15:0] flash_cfg_reg_rddata    ,

output wire        SLAVE_CLK               , //向AXI总线提供的本主机时钟信号
output wire        SLAVE_RSTN              , //向AXI总线提供的本主机复位信号
input  wire [ 3:0] SLAVE_WR_ADDR_ID        , //写地址通道-ID
input  wire [31:0] SLAVE_WR_ADDR           , //写地址通道-地址
input  wire [ 7:0] SLAVE_WR_ADDR_LEN       , //写地址通道-突发长度-最小为0（1突发），最大为255（256突发）
input  wire [ 1:0] SLAVE_WR_ADDR_BURST     , //写地址通道-突发类型
input  wire        SLAVE_WR_ADDR_VALID     , //写地址通道-握手信号-有效
output reg         SLAVE_WR_ADDR_READY     , //写地址通道-握手信号-准备
input  wire [31:0] SLAVE_WR_DATA           , //写数据通道-数据
input  wire [ 3:0] SLAVE_WR_STRB           , //写数据通道-选通
input  wire        SLAVE_WR_DATA_LAST      , //写数据通道-last信号
input  wire        SLAVE_WR_DATA_VALID     , //写数据通道-握手信号-有效
output reg         SLAVE_WR_DATA_READY     , //写数据通道-握手信号-准备
output reg  [ 3:0] SLAVE_WR_BACK_ID        , //写响应通道-ID
output reg  [ 1:0] SLAVE_WR_BACK_RESP      , //写响应通道-响应 //SLAVE_WR_DATA_LAST拉高的同时或者之后 00 01正常 10写错误 11地址有问题找不到从机
output reg         SLAVE_WR_BACK_VALID     , //写响应通道-握手信号-有效
input  wire        SLAVE_WR_BACK_READY     , //写响应通道-握手信号-准备
input  wire [ 3:0] SLAVE_RD_ADDR_ID        , //读地址通道-ID
input  wire [31:0] SLAVE_RD_ADDR           , //读地址通道-地址
input  wire [ 7:0] SLAVE_RD_ADDR_LEN       , //读地址通道-突发长度。最小为0（1突发），最大为255（256突发）
input  wire [ 1:0] SLAVE_RD_ADDR_BURST     , //读地址通道-突发类型。
input  wire        SLAVE_RD_ADDR_VALID     , //读地址通道-握手信号-有效
output reg         SLAVE_RD_ADDR_READY     , //读地址通道-握手信号-准备
output reg  [ 3:0] SLAVE_RD_BACK_ID        , //读数据通道-ID
output reg  [31:0] SLAVE_RD_DATA           , //读数据通道-数据
output reg  [ 1:0] SLAVE_RD_DATA_RESP      , //读数据通道-响应
output reg         SLAVE_RD_DATA_LAST      , //读数据通道-last信号
output reg         SLAVE_RD_DATA_VALID     , //读数据通道-握手信号-有效
input  wire        SLAVE_RD_DATA_READY       //读数据通道-握手信号-准备
);

//读/写FLASH芯片配置寄存器及状态指示信号
assign flash_cfg_cmd_en     = 0;
assign flash_cfg_cmd        = 0;
assign flash_cfg_reg_wrdata = 0;

/*
ADDR: 0X00: 写Flash-读写地址——控制位
[31:16]: wr_sector_num
[15: 0]: {flash_wr_en,-,-,-, start_wr_sector}

ADDR: 0X01: 写Flash-只写地址——FIFO入口
[31:0]:  写比特流数据入口

ADDR: 0X02: 写Flash-只读地址——标志位
[31:24]: {-, -, -, -, -, -, -,      wr_fifo_full}
[23:16]: {-, -, -, -, -, -, -,     wr_fifo_empty}
[15: 8]: {-, -, -, -, -, -, -,     flash_wr_done}
[ 7: 0]: {-, -, -, -, -, -, -,  flash_clear_done}

ADDR: 0X03: 读Flash-读写地址——控制位1
[31:16]: rd_sector_num
[15: 0]: {flash_rd_en,-,-,-, start_rd_sub_sector}

ADDR: 0X04: 读Flash-读写地址——控制位2
[31:24]: {                                            }
[23:16]: {-, -, -, -, -, -,{   bs_crc32_ok           }}
[15: 8]: {-, -, -, -, -, -, -,            crc_check_en}
[ 7: 0]: {-, -, -, -, -, -, -,     bitstream_up2cpu_en}

ADDR: 0X05: 读Flash-只读地址——FIFO出口
[31:0]: 读比特流数据出口

ADDR: 0X06: 读Flash-只读地址——CRC校验值
[31:0]: CRC校验值 bs_readback_crc

ADDR: 0X07: 读Flash-只读地址——标志位
[31:24]: {-, -, -, -, -, -, -,         rd_fifo_afull}
[23:16]: {-, -, -, -, -, -, -,         rd_fifo_empty}
[15: 8]: {-, -, -, -, -, -, -,         flash_rd_done}
[ 7: 0]: {-, -, -, -, -, -, -, bs_readback_crc_valid}

ADDR: 0X08: 热启动开关-读写地址——控制位
[31: 8]: hotreset_addr
[ 7: 0]: {-, -, -, -, -, -, -,    hotreset_en}

ADDR: 0X09: 只读地址 版本号
[31: 0]: FPGA_VERSION[31:0]
*/

localparam RU_WRBIT_RW_CTRL_ADDR = 32'h0000_0000;
localparam RU_WRBIT_WO_FIFO_ADDR = 32'h0000_0001;
localparam RU_WRBIT_RO_FLAG_ADDR = 32'h0000_0002;
  
localparam RU_RDBIT_RW_CTRL1_ADDR = 32'h0000_0003;
localparam RU_RDBIT_RW_CTRL2_ADDR = 32'h0000_0004;
localparam RU_RDBIT_RO_FIFO_ADDR = 32'h0000_0005;
localparam RU_RDBIT_RO__CRC_ADDR = 32'h0000_0006;
localparam RU_RDBIT_RO_FLAG_ADDR = 32'h0000_0007;
  
localparam RU_HOTRS_RW_CTRL_ADDR = 32'h0000_0008;
localparam RU_FPGAV_RO_ADDR      = 32'h0000_0009;

assign SLAVE_CLK = clk;
wire SLAVE_RSTN_SYNC;
rstn_sync ru_rstn_sync(clk,rstn,SLAVE_RSTN_SYNC);
assign SLAVE_RSTN = SLAVE_RSTN_SYNC;

reg  [ 3:0] wr_addr_id;   
reg  [31:0] wr_addr;
reg  [ 1:0] wr_addr_burst;
reg         wr_error_detect;
reg  [ 1:0] cu_wr_st, nt_wr_st;
localparam ST_WR_IDLE = 2'b00,
           ST_WR_DATA = 2'b01,
           ST_WR_RESP = 2'b10;

reg  [ 3:0] rd_addr_id;   
reg  [31:0] rd_addr;
reg  [ 7:0] rd_addr_len;
reg  [ 1:0] rd_addr_burst;
reg         rd_error_detect, rd_error_detect_reg;
reg  [ 7:0] trans_num;
reg         cu_rd_st, nt_rd_st;
localparam ST_RD_IDLE = 1'b0,
           ST_RD_DATA = 1'b1;

wire        wr_fifo_rst;
wire        wr_fifo_wr_en;
wire [31:0] wr_fifo_wr_data;
wire        wr_fifo_rd_en;
wire [ 7:0] wr_fifo_rd_data;
reg         wr_fifo_rd_data_valid;
wire        wr_fifo_full;
wire        wr_fifo_empty;
wire [11:0] wr_fifo_bytes_num;
reg  [11:0] wr_fifo_trans_cnt;

wire        rd_fifo_rst;
wire        rd_fifo_wr_en;
wire [ 7:0] rd_fifo_wr_data;
wire        rd_fifo_rd_en;
wire [31:0] rd_fifo_rd_data;
reg         rd_fifo_rd_data_valid;
wire        rd_fifo_afull;
wire        rd_fifo_empty;

//___________________写通道___________________//

always @(*) begin
    if(~SLAVE_RSTN_SYNC) nt_wr_st <= ST_WR_IDLE;
    else case (cu_wr_st)
        ST_WR_IDLE: nt_wr_st <= (SLAVE_WR_ADDR_READY && SLAVE_WR_ADDR_VALID)?(ST_WR_DATA):(ST_WR_IDLE);
        ST_WR_DATA: nt_wr_st <= (SLAVE_WR_DATA_READY && SLAVE_WR_DATA_VALID && SLAVE_WR_DATA_LAST)?(ST_WR_RESP):(ST_WR_DATA);
        ST_WR_RESP: nt_wr_st <= (SLAVE_WR_BACK_READY && SLAVE_WR_BACK_VALID)?(ST_WR_IDLE):(ST_WR_RESP);
        default:    nt_wr_st <= ST_WR_IDLE;
    endcase
end
always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) cu_wr_st <= ST_WR_IDLE;
    else cu_wr_st <= nt_wr_st;
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) begin
        wr_addr_id <= 0;
        wr_addr_burst <= 0;
    end else if(SLAVE_WR_ADDR_READY && SLAVE_WR_ADDR_VALID)begin
        wr_addr_id <= SLAVE_WR_ADDR_ID;
        wr_addr_burst <= SLAVE_WR_ADDR_BURST;
    end else begin
        wr_addr_id <= wr_addr_id;
        wr_addr_burst <= wr_addr_burst;
    end
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) wr_addr <= 0;
    else if(SLAVE_WR_ADDR_READY && SLAVE_WR_ADDR_VALID) wr_addr <= SLAVE_WR_ADDR - OFFSET_ADDR;
    else if((cu_wr_st == ST_WR_DATA) && SLAVE_WR_DATA_READY && SLAVE_WR_DATA_VALID && (wr_addr_burst == 2'b01)) wr_addr <= wr_addr + 1;
    else wr_addr <= wr_addr;
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) wr_error_detect <= 0;
    else if(cu_wr_st == ST_WR_IDLE) wr_error_detect <= 0;
    else if(cu_wr_st == ST_WR_DATA)begin
        if((wr_addr_burst == 2'b10) || (wr_addr_burst == 2'b11)) wr_error_detect <= 1;
        else if((wr_addr < RU_WRBIT_RW_CTRL_ADDR) || (wr_addr > RU_FPGAV_RO_ADDR)) wr_error_detect <= 1;
        else if((wr_addr == RU_WRBIT_RO_FLAG_ADDR) ||
                (wr_addr == RU_RDBIT_RO_FIFO_ADDR) ||
                (wr_addr == RU_RDBIT_RO_FLAG_ADDR) ||
                (wr_addr == RU_RDBIT_RO__CRC_ADDR) ||
                (wr_addr == RU_FPGAV_RO_ADDR)) wr_error_detect <= 1;
        else wr_error_detect <= 0;
    end else wr_error_detect <= wr_error_detect;
end

assign SLAVE_WR_ADDR_READY = (cu_wr_st == ST_WR_IDLE);
assign SLAVE_WR_BACK_ID    = wr_addr_id;
assign SLAVE_WR_BACK_RESP  = (wr_error_detect)?(2'b10):(2'b00);
assign SLAVE_WR_BACK_VALID = (cu_wr_st == ST_WR_RESP);

//___________________读通道___________________//

// always @(posedge clk) begin
//     if(~SLAVE_RSTN_SYNC) led <= 0;
//     else if(SLAVE_WR_DATA_READY && SLAVE_WR_DATA_VALID && (wr_addr == ADDR))begin
//         led <= SLAVE_WR_DATA;
//         $display("%m: at time %0t INFO: remote update slave recv write data %h", $time, SLAVE_WR_DATA);
//     end else led <= led;
// end

always @(*) begin
    if(~SLAVE_RSTN_SYNC) nt_rd_st <= ST_RD_IDLE;
    else case (cu_rd_st)
        ST_RD_IDLE: nt_rd_st <= (SLAVE_RD_ADDR_READY && SLAVE_RD_ADDR_VALID)?(ST_RD_DATA):(ST_RD_IDLE);
        ST_RD_DATA: nt_rd_st <= (SLAVE_RD_DATA_READY && SLAVE_RD_DATA_VALID && SLAVE_RD_DATA_LAST)?(ST_RD_IDLE):(ST_RD_DATA);
    endcase
end
always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) cu_rd_st <= ST_RD_IDLE;
    else cu_rd_st <= nt_rd_st;
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) begin
        rd_addr_id <= 0;
        rd_addr_burst <= 0;
        rd_addr_len <= 0;
    end else if(SLAVE_RD_ADDR_READY && SLAVE_RD_ADDR_VALID)begin
        rd_addr_id <= SLAVE_RD_ADDR_ID;
        rd_addr_burst <= SLAVE_RD_ADDR_BURST;
        rd_addr_len <= SLAVE_RD_ADDR_LEN;
    end else begin
        rd_addr_id <= rd_addr_id;
        rd_addr_burst <= rd_addr_burst;
        rd_addr_len <= rd_addr_len;
    end
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) rd_addr <= 0;
    else if(SLAVE_RD_ADDR_READY && SLAVE_RD_ADDR_VALID) rd_addr <= SLAVE_RD_ADDR - OFFSET_ADDR;
    else if((cu_rd_st == ST_RD_DATA) && SLAVE_RD_DATA_READY && SLAVE_RD_DATA_VALID && (rd_addr_burst == 2'b01)) rd_addr <= rd_addr + 1;
    else rd_addr <= rd_addr;
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) trans_num <= 0;
    else if(cu_rd_st == ST_RD_IDLE) trans_num <= 0;
    else if(SLAVE_RD_DATA_READY && SLAVE_RD_DATA_VALID) trans_num <= trans_num + 1;
    else trans_num <= trans_num;
end

always @(*) begin
    if(~SLAVE_RSTN_SYNC) rd_error_detect <= 0;
    else if(cu_rd_st == ST_RD_DATA)begin
        if((rd_addr_burst == 2'b10) || (rd_addr_burst == 2'b11)) rd_error_detect <= 1;
        if((rd_addr < RU_WRBIT_RW_CTRL_ADDR) || (rd_addr > RU_FPGAV_RO_ADDR)) rd_error_detect <= 1;
        else if(rd_addr == RU_WRBIT_WO_FIFO_ADDR) rd_error_detect <= 1;
        else rd_error_detect <= 0;
    end else rd_error_detect <= 0;
end
always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) rd_error_detect_reg <= 0;
    else rd_error_detect_reg <= rd_error_detect;
end

assign SLAVE_RD_ADDR_READY = (cu_rd_st == ST_RD_IDLE);
assign SLAVE_RD_BACK_ID    = rd_addr_id;
assign SLAVE_RD_DATA_RESP  = (rd_error_detect || rd_error_detect_reg)?(2'b10):(2'b00);
assign SLAVE_RD_DATA_LAST  = (SLAVE_RD_DATA_VALID && (trans_num == rd_addr_len));

//写通道的READY信号
always @(*) begin
    if(~SLAVE_RSTN_SYNC || (cu_wr_st == ST_WR_IDLE) || (cu_wr_st == ST_WR_RESP)) SLAVE_WR_DATA_READY <= 0;
    else if(cu_wr_st == ST_WR_DATA)begin
        case (wr_addr)
            RU_WRBIT_WO_FIFO_ADDR: SLAVE_WR_DATA_READY <= (~wr_fifo_full);
            default                   : SLAVE_WR_DATA_READY <= 1;
        endcase
    end else SLAVE_WR_DATA_READY <= 0;
end

//读通道的VALID信号
always @(*) begin
    if(~SLAVE_RSTN_SYNC || (cu_rd_st == ST_RD_IDLE)) SLAVE_RD_DATA_VALID <= 0;
    else if(cu_rd_st == ST_RD_DATA)begin
        case (rd_addr)
            RU_RDBIT_RO_FIFO_ADDR: SLAVE_RD_DATA_VALID <= (rd_fifo_rd_data_valid);
            default                   : SLAVE_RD_DATA_VALID <= 1;
        endcase
    end else SLAVE_RD_DATA_VALID <= 0;
end

//读通道的DATA选通
always @(*) begin
    if(~SLAVE_RSTN_SYNC || (cu_rd_st == ST_RD_IDLE)) SLAVE_RD_DATA <= 0;
    else if(cu_rd_st == ST_RD_DATA)begin
        case (rd_addr)
            RU_WRBIT_RW_CTRL_ADDR: SLAVE_RD_DATA <= {wr_sector_num[15:0],flash_wr_en,3'b0,start_wr_sector[11:0]};
            RU_WRBIT_WO_FIFO_ADDR: SLAVE_RD_DATA <= 32'hFFFF_FFFF;
            RU_WRBIT_RO_FLAG_ADDR: SLAVE_RD_DATA <= {{7'b0,wr_fifo_full},{7'b0,wr_fifo_empty},{7'b0,flash_wr_done},{7'b0, flash_clear_done}};
            RU_RDBIT_RW_CTRL1_ADDR:SLAVE_RD_DATA <= {rd_sector_num[15:0],flash_rd_en,3'b0,start_rd_sub_sector[11:0]};
            RU_RDBIT_RW_CTRL2_ADDR:SLAVE_RD_DATA <= {{8'b0},{6'b0,bs_crc32_ok},{7'b0,crc_check_en} ,{7'b0, bitstream_up2cpu_en}};
            RU_RDBIT_RO_FIFO_ADDR: SLAVE_RD_DATA <= rd_fifo_rd_data;
            RU_RDBIT_RO__CRC_ADDR: SLAVE_RD_DATA <= bs_readback_crc;
            RU_RDBIT_RO_FLAG_ADDR: SLAVE_RD_DATA <= {{7'b0,rd_fifo_afull},{7'b0,rd_fifo_empty},{7'b0,flash_rd_done},{7'b0, bs_readback_crc_valid}};
            RU_HOTRS_RW_CTRL_ADDR: SLAVE_RD_DATA <= {hotreset_addr,{7'b0, hotreset_en}};
            RU_FPGAV_RO_ADDR     : SLAVE_RD_DATA <= FPGA_VERSION[31:0];
            default              : SLAVE_RD_DATA <= 32'hFFFF_FFFF;
        endcase
    end else SLAVE_RD_DATA <= 32'hFFFF_FFFF;
end

assign wr_fifo_rst     = (~SLAVE_RSTN_SYNC);
assign wr_fifo_wr_en   = (cu_wr_st == ST_WR_DATA) && (wr_addr == RU_WRBIT_WO_FIFO_ADDR) && (SLAVE_WR_DATA_VALID) && (SLAVE_WR_DATA_READY);
assign wr_fifo_wr_data = SLAVE_WR_DATA;
assign wr_fifo_rd_en   = (~wr_fifo_empty) && ((~wr_fifo_rd_data_valid) || (bitstream_valid));
always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) wr_fifo_rd_data_valid <= 0;
    else if((~wr_fifo_rd_data_valid) && (~wr_fifo_empty) && (wr_fifo_rd_en)) wr_fifo_rd_data_valid <= 1;
    else if((wr_fifo_rd_data_valid) && (wr_fifo_empty) && (bitstream_valid)) wr_fifo_rd_data_valid <= 0;
    else wr_fifo_rd_data_valid <= wr_fifo_rd_data_valid;
end

assign rd_fifo_rst     = (~SLAVE_RSTN_SYNC);
assign rd_fifo_wr_en   = flash_rd_valid;
assign rd_fifo_wr_data = flash_rd_data;
assign rd_fifo_rd_en   = (~rd_fifo_empty) && ((~rd_fifo_rd_data_valid) || ((cu_rd_st == ST_RD_DATA) && (rd_addr == RU_RDBIT_RO_FIFO_ADDR) && (SLAVE_RD_DATA_VALID) && (SLAVE_RD_DATA_READY)));
always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) rd_fifo_rd_data_valid <= 0;
    else if((~rd_fifo_rd_data_valid) && (~rd_fifo_empty) && (rd_fifo_rd_en)) rd_fifo_rd_data_valid <= 1;
    else if((rd_fifo_rd_data_valid) && (rd_fifo_empty) && ((cu_rd_st == ST_RD_DATA) && (rd_addr == RU_RDBIT_RO_FIFO_ADDR) && (SLAVE_RD_DATA_VALID) && (SLAVE_RD_DATA_READY)))
        rd_fifo_rd_data_valid <= 0;
    else rd_fifo_rd_data_valid <= rd_fifo_rd_data_valid;
end


reg cu_wr_fifo_st, nt_wr_fifo_st;
localparam ST_WR_FIFO_IDLE  = 1'b0;
localparam ST_WR_FIFO_TRANS = 1'b1;
always @(*) begin
    if(~SLAVE_RSTN_SYNC) nt_wr_fifo_st <= ST_WR_FIFO_IDLE;
    else case(cu_wr_fifo_st)
        ST_WR_FIFO_IDLE : nt_wr_fifo_st <= (wr_fifo_bytes_num >= 255)?(ST_WR_FIFO_TRANS):(ST_WR_FIFO_IDLE); //因为会事先读出来一个
        ST_WR_FIFO_TRANS: nt_wr_fifo_st <= (bitstream_eop && bitstream_valid)?(ST_WR_FIFO_IDLE):(ST_WR_FIFO_TRANS);
    endcase
end
always @(posedge clk or negedge SLAVE_RSTN_SYNC)begin
    if(~SLAVE_RSTN_SYNC) cu_wr_fifo_st <= ST_WR_FIFO_IDLE;
    else cu_wr_fifo_st <= nt_wr_fifo_st;
end  

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC) wr_fifo_trans_cnt <= 0;
    else if(cu_wr_fifo_st == ST_WR_FIFO_TRANS) begin
        if(bitstream_valid) wr_fifo_trans_cnt <= wr_fifo_trans_cnt + 1;
        else wr_fifo_trans_cnt <= wr_fifo_trans_cnt;
    end else wr_fifo_trans_cnt <= 0;
end
assign bitstream_fifo_rd_rdy = (cu_wr_fifo_st == ST_WR_FIFO_TRANS);
assign bitstream_valid = bitstream_fifo_rd_req;
assign bitstream_data = wr_fifo_rd_data;
assign bitstream_eop = (wr_fifo_trans_cnt >= 255) & bitstream_valid;
assign flash_rd_data_fifo_afull = rd_fifo_afull;

remote_update_wr_fifo remote_update_wr_fifo_inst(
    .clk           (clk),
    .rst           (wr_fifo_rst),
    .wr_en         (wr_fifo_wr_en),
    .wr_data       (wr_fifo_wr_data),
    .rd_en         (wr_fifo_rd_en),
    .rd_data       (wr_fifo_rd_data),

    .wr_full       (wr_fifo_full),
    .rd_empty      (wr_fifo_empty),
    .rd_water_level(wr_fifo_bytes_num)
);

remote_update_rd_fifo remote_update_rd_fifo_inst(
    .clk           (clk),
    .rst           (rd_fifo_rst),
    .wr_en         (rd_fifo_wr_en),
    .wr_data       (rd_fifo_wr_data),
    .rd_en         (rd_fifo_rd_en),
    .rd_data       (rd_fifo_rd_data),

    .rd_empty      (rd_fifo_empty),
    .almost_full   (rd_fifo_afull) //set n-256 bytes almost full
);

///__________输出信号___________///
always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC)begin
        flash_wr_en <= 0;
        start_wr_sector <= 0;
        wr_sector_num <= 0;
    end else if(SLAVE_WR_DATA_VALID && SLAVE_WR_DATA_READY && wr_addr == RU_WRBIT_RW_CTRL_ADDR)begin
        wr_sector_num[15:8]       <= (SLAVE_WR_STRB[3])?(SLAVE_WR_DATA[31:24]):(wr_sector_num[15:8]      );
        wr_sector_num[ 7:0]       <= (SLAVE_WR_STRB[2])?(SLAVE_WR_DATA[23:16]):(wr_sector_num[ 7:0]      );
        flash_wr_en               <= (SLAVE_WR_STRB[1])?(SLAVE_WR_DATA[   15]):(flash_wr_en              );
        start_wr_sector[11:8] <= (SLAVE_WR_STRB[1])?(SLAVE_WR_DATA[11: 8]):(start_wr_sector[11:8]);
        start_wr_sector[ 7:0] <= (SLAVE_WR_STRB[0])?(SLAVE_WR_DATA[ 7: 0]):(start_wr_sector[ 7:0]);
    end else begin
        flash_wr_en <= 0;
        start_wr_sector <= start_wr_sector;
        wr_sector_num <= wr_sector_num;
    end
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC)begin
        flash_rd_en <= 0;
        start_rd_sub_sector <= 0;
        rd_sector_num <= 0;
    end else if(SLAVE_WR_DATA_VALID && SLAVE_WR_DATA_READY && wr_addr == RU_RDBIT_RW_CTRL1_ADDR)begin
        rd_sector_num[15:8]       <= (SLAVE_WR_STRB[3])?(SLAVE_WR_DATA[31:24]):(rd_sector_num[15:8]      );
        rd_sector_num[ 7:0]       <= (SLAVE_WR_STRB[2])?(SLAVE_WR_DATA[23:16]):(rd_sector_num[ 7:0]      );
        flash_rd_en               <= (SLAVE_WR_STRB[1])?(SLAVE_WR_DATA[   15]):(flash_rd_en              );
        start_rd_sub_sector[11:8] <= (SLAVE_WR_STRB[1])?(SLAVE_WR_DATA[11: 8]):(start_rd_sub_sector[11:8]);
        start_rd_sub_sector[ 7:0] <= (SLAVE_WR_STRB[0])?(SLAVE_WR_DATA[ 7: 0]):(start_rd_sub_sector[ 7:0]);
    end else begin
        flash_rd_en <= 0;
        start_rd_sub_sector <= start_rd_sub_sector;
        rd_sector_num <= rd_sector_num;
    end
end

always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC)begin
        bs_crc32_ok                      <= 0;
        crc_check_en                     <= 0;
        bitstream_up2cpu_en              <= 0;
    end else if(SLAVE_WR_DATA_VALID && SLAVE_WR_DATA_READY && wr_addr == RU_RDBIT_RW_CTRL2_ADDR)begin
        bs_crc32_ok                      <= (SLAVE_WR_STRB[2])?(SLAVE_WR_DATA[17:16]):(bs_crc32_ok        );
        crc_check_en                     <= (SLAVE_WR_STRB[1])?(SLAVE_WR_DATA[8]    ):(crc_check_en       );
        bitstream_up2cpu_en              <= (SLAVE_WR_STRB[0])?(SLAVE_WR_DATA[0]    ):(bitstream_up2cpu_en);
    end else begin
        bs_crc32_ok                      <= bs_crc32_ok                     ;
        crc_check_en                     <= crc_check_en                    ;
        bitstream_up2cpu_en              <= bitstream_up2cpu_en             ;
    end
end
always @(posedge clk or negedge SLAVE_RSTN_SYNC) begin
    if(~SLAVE_RSTN_SYNC)begin
        hotreset_addr <= 0;
        hotreset_en <= 0;
    end else if(SLAVE_WR_DATA_VALID && SLAVE_WR_DATA_READY && wr_addr == RU_HOTRS_RW_CTRL_ADDR)begin
        hotreset_addr[23:16] <= (SLAVE_WR_STRB[3])?(SLAVE_WR_DATA[31:24]):(hotreset_addr[23:16]);
        hotreset_addr[15: 8] <= (SLAVE_WR_STRB[2])?(SLAVE_WR_DATA[23:16]):(hotreset_addr[15: 8]);
        hotreset_addr[ 7: 0] <= (SLAVE_WR_STRB[1])?(SLAVE_WR_DATA[15: 8]):(hotreset_addr[ 7: 0]);
        hotreset_en   <= (SLAVE_WR_STRB[0])?(SLAVE_WR_DATA[0]):(hotreset_en);
    end else begin
        hotreset_addr <= hotreset_addr;
        hotreset_en <= 0;//自动置0
    end
end

endmodule