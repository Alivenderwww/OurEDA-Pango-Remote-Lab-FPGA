module decoder_5_32 (
    input [4:0] in,
    output reg [31:0] sel
);
    always@(*)begin
        case(in)
            5'd0  : sel = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            5'd1  : sel = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            5'd2  : sel = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
            5'd3  : sel = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
            5'd4  : sel = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
            5'd5  : sel = 32'b0000_0000_0000_0000_0000_0000_0010_0000;
            5'd6  : sel = 32'b0000_0000_0000_0000_0000_0000_0100_0000;
            5'd7  : sel = 32'b0000_0000_0000_0000_0000_0000_1000_0000;
            5'd8  : sel = 32'b0000_0000_0000_0000_0000_0001_0000_0000;
            5'd9  : sel = 32'b0000_0000_0000_0000_0000_0010_0000_0000;
            5'd10 : sel = 32'b0000_0000_0000_0000_0000_0100_0000_0000;
            5'd11 : sel = 32'b0000_0000_0000_0000_0000_1000_0000_0000;
            5'd12 : sel = 32'b0000_0000_0000_0000_0001_0000_0000_0000;
            5'd13 : sel = 32'b0000_0000_0000_0000_0010_0000_0000_0000;
            5'd14 : sel = 32'b0000_0000_0000_0000_0100_0000_0000_0000;
            5'd15 : sel = 32'b0000_0000_0000_0000_1000_0000_0000_0000;
            5'd16 : sel = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
            5'd17 : sel = 32'b0000_0000_0000_0010_0000_0000_0000_0000;
            5'd18 : sel = 32'b0000_0000_0000_0100_0000_0000_0000_0000;
            5'd19 : sel = 32'b0000_0000_0000_1000_0000_0000_0000_0000;
            5'd20 : sel = 32'b0000_0000_0001_0000_0000_0000_0000_0000;
            5'd21 : sel = 32'b0000_0000_0010_0000_0000_0000_0000_0000;
            5'd22 : sel = 32'b0000_0000_0100_0000_0000_0000_0000_0000;
            5'd23 : sel = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
            5'd24 : sel = 32'b0000_0001_0000_0000_0000_0000_0000_0000;
            5'd25 : sel = 32'b0000_0010_0000_0000_0000_0000_0000_0000;
            5'd26 : sel = 32'b0000_0100_0000_0000_0000_0000_0000_0000;
            5'd27 : sel = 32'b0000_1000_0000_0000_0000_0000_0000_0000;
            5'd28 : sel = 32'b0001_0000_0000_0000_0000_0000_0000_0000;
            5'd29 : sel = 32'b0010_0000_0000_0000_0000_0000_0000_0000;
            5'd30 : sel = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
            5'd31 : sel = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
        endcase
    end
endmodule